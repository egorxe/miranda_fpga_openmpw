VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1426.380 2924.800 1427.580 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3486.100 2.400 3487.300 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3224.980 2.400 3226.180 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2964.540 2.400 2965.740 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1692.260 2924.800 1693.460 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2703.420 2.400 2704.620 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2442.980 2.400 2444.180 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2182.540 2.400 2183.740 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1921.420 2.400 1922.620 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1660.980 2.400 1662.180 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1399.860 2.400 1401.060 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1139.420 2.400 1140.620 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 878.980 2.400 880.180 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 617.860 2.400 619.060 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1958.140 2924.800 1959.340 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2223.340 2924.800 2224.540 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2489.220 2924.800 2490.420 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2755.100 2924.800 2756.300 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3020.300 2924.800 3021.500 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3286.180 2924.800 3287.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 32.380 2924.800 33.580 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2289.980 2924.800 2291.180 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2555.860 2924.800 2557.060 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2821.060 2924.800 2822.260 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3086.940 2924.800 3088.140 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3352.820 2924.800 3354.020 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 230.940 2924.800 232.140 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3420.820 2.400 3422.020 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3159.700 2.400 3160.900 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2899.260 2.400 2900.460 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2638.820 2.400 2640.020 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2377.700 2.400 2378.900 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2117.260 2.400 2118.460 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 430.180 2924.800 431.380 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1856.140 2.400 1857.340 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1595.700 2.400 1596.900 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1335.260 2.400 1336.460 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1074.140 2.400 1075.340 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 813.700 2.400 814.900 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 552.580 2.400 553.780 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 357.420 2.400 358.620 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 161.580 2.400 162.780 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 629.420 2924.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 828.660 2924.800 829.860 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1027.900 2924.800 1029.100 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1227.140 2924.800 1228.340 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1493.020 2924.800 1494.220 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1758.900 2924.800 1760.100 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2024.100 2924.800 2025.300 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 164.980 2924.800 166.180 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2422.580 2924.800 2423.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2688.460 2924.800 2689.660 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2954.340 2924.800 2955.540 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3219.540 2924.800 3220.740 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3485.420 2924.800 3486.620 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 364.220 2924.800 365.420 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3290.260 2.400 3291.460 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3029.820 2.400 3031.020 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.700 2.400 2769.900 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2508.260 2.400 2509.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2247.140 2.400 2248.340 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1986.700 2.400 1987.900 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 563.460 2924.800 564.660 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1726.260 2.400 1727.460 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1465.140 2.400 1466.340 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 2.400 1205.900 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 943.580 2.400 944.780 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 683.140 2.400 684.340 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 422.700 2.400 423.900 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 226.860 2.400 228.060 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 31.700 2.400 32.900 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 762.700 2924.800 763.900 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 961.940 2924.800 963.140 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1161.180 2924.800 1162.380 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1360.420 2924.800 1361.620 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1625.620 2924.800 1626.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1891.500 2924.800 1892.700 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2157.380 2924.800 2158.580 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 98.340 2924.800 99.540 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2356.620 2924.800 2357.820 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2621.820 2924.800 2623.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2887.700 2924.800 2888.900 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3153.580 2924.800 3154.780 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3418.780 2924.800 3419.980 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 297.580 2924.800 298.780 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3355.540 2.400 3356.740 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3095.100 2.400 3096.300 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2833.980 2.400 2835.180 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2573.540 2.400 2574.740 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2312.420 2.400 2313.620 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2051.980 2.400 2053.180 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 496.820 2924.800 498.020 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1791.540 2.400 1792.740 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1530.420 2.400 1531.620 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1269.980 2.400 1271.180 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1008.860 2.400 1010.060 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 2.400 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 487.300 2.400 488.500 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 292.140 2.400 293.340 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 96.300 2.400 97.500 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 696.060 2924.800 697.260 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 895.300 2924.800 896.500 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1094.540 2924.800 1095.740 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1293.780 2924.800 1294.980 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1559.660 2924.800 1560.860 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1824.860 2924.800 1826.060 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2090.740 2924.800 2091.940 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 629.230 -4.800 629.790 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.530 -4.800 2403.090 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2420.010 -4.800 2420.570 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2437.950 -4.800 2438.510 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2473.370 -4.800 2473.930 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2490.850 -4.800 2491.410 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2508.790 -4.800 2509.350 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2526.730 -4.800 2527.290 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2544.210 -4.800 2544.770 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2562.150 -4.800 2562.710 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.330 -4.800 806.890 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2597.570 -4.800 2598.130 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.050 -4.800 2615.610 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.990 -4.800 2633.550 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2650.470 -4.800 2651.030 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2668.410 -4.800 2668.970 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2685.890 -4.800 2686.450 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2721.770 -4.800 2722.330 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.250 -4.800 2739.810 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2757.190 -4.800 2757.750 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2774.670 -4.800 2775.230 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.610 -4.800 2793.170 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2810.090 -4.800 2810.650 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2828.030 -4.800 2828.590 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2845.510 -4.800 2846.070 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2863.450 -4.800 2864.010 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2881.390 -4.800 2881.950 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 841.750 -4.800 842.310 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 859.690 -4.800 860.250 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 877.170 -4.800 877.730 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 895.110 -4.800 895.670 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 930.530 -4.800 931.090 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 646.710 -4.800 647.270 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.370 -4.800 1001.930 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1054.730 -4.800 1055.290 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.210 -4.800 1072.770 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1090.150 -4.800 1090.710 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1107.630 -4.800 1108.190 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.570 -4.800 1126.130 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1143.510 -4.800 1144.070 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.650 -4.800 665.210 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1178.930 -4.800 1179.490 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.410 -4.800 1196.970 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1214.350 -4.800 1214.910 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1231.830 -4.800 1232.390 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.770 -4.800 1250.330 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1267.250 -4.800 1267.810 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1303.130 -4.800 1303.690 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.610 -4.800 1321.170 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 682.130 -4.800 682.690 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1338.550 -4.800 1339.110 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.030 -4.800 1356.590 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.970 -4.800 1374.530 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1391.450 -4.800 1392.010 2.400 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1426.870 -4.800 1427.430 2.400 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1444.810 -4.800 1445.370 2.400 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1462.750 -4.800 1463.310 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1480.230 -4.800 1480.790 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1498.170 -4.800 1498.730 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1515.650 -4.800 1516.210 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1551.070 -4.800 1551.630 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.010 -4.800 1569.570 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.490 -4.800 1587.050 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1604.430 -4.800 1604.990 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1639.850 -4.800 1640.410 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1675.270 -4.800 1675.830 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 717.550 -4.800 718.110 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.210 -4.800 1693.770 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.690 -4.800 1711.250 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1728.630 -4.800 1729.190 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1764.050 -4.800 1764.610 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.530 -4.800 1782.090 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1799.470 -4.800 1800.030 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.410 -4.800 1817.970 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.890 -4.800 1835.450 2.400 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1852.830 -4.800 1853.390 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.490 -4.800 736.050 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1888.250 -4.800 1888.810 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1923.670 -4.800 1924.230 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1976.570 -4.800 1977.130 2.400 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2029.930 -4.800 2030.490 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.970 -4.800 753.530 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2047.870 -4.800 2048.430 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2065.350 -4.800 2065.910 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2083.290 -4.800 2083.850 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2100.770 -4.800 2101.330 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2136.190 -4.800 2136.750 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.130 -4.800 2154.690 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2172.070 -4.800 2172.630 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2189.550 -4.800 2190.110 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.490 -4.800 2208.050 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 770.910 -4.800 771.470 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2224.970 -4.800 2225.530 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2260.390 -4.800 2260.950 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.330 -4.800 2278.890 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.810 -4.800 2296.370 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2313.750 -4.800 2314.310 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2349.170 -4.800 2349.730 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2384.590 -4.800 2385.150 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.850 -4.800 789.410 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 634.750 -4.800 635.310 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.990 -4.800 2426.550 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2443.930 -4.800 2444.490 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2461.410 -4.800 2461.970 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2479.350 -4.800 2479.910 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2514.770 -4.800 2515.330 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.250 -4.800 2532.810 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2550.190 -4.800 2550.750 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2567.670 -4.800 2568.230 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 812.310 -4.800 812.870 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.610 -4.800 2586.170 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2603.550 -4.800 2604.110 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 2.400 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2638.970 -4.800 2639.530 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.450 -4.800 2657.010 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2674.390 -4.800 2674.950 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2691.870 -4.800 2692.430 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.810 -4.800 2710.370 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2727.290 -4.800 2727.850 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 830.250 -4.800 830.810 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2763.170 -4.800 2763.730 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2780.650 -4.800 2781.210 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2798.590 -4.800 2799.150 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2816.070 -4.800 2816.630 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2834.010 -4.800 2834.570 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2851.490 -4.800 2852.050 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2869.430 -4.800 2869.990 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 847.730 -4.800 848.290 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 883.150 -4.800 883.710 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.090 -4.800 901.650 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 936.510 -4.800 937.070 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.690 -4.800 653.250 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.410 -4.800 989.970 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.770 -4.800 1043.330 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1060.710 -4.800 1061.270 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1096.130 -4.800 1096.690 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1113.610 -4.800 1114.170 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1131.550 -4.800 1132.110 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.030 -4.800 1149.590 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 670.630 -4.800 671.190 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.970 -4.800 1167.530 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1184.910 -4.800 1185.470 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 2.400 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1220.330 -4.800 1220.890 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1237.810 -4.800 1238.370 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1255.750 -4.800 1256.310 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1273.230 -4.800 1273.790 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1291.170 -4.800 1291.730 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1308.650 -4.800 1309.210 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 688.110 -4.800 688.670 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1344.070 -4.800 1344.630 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.010 -4.800 1362.570 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.950 -4.800 1380.510 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1397.430 -4.800 1397.990 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1415.370 -4.800 1415.930 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1432.850 -4.800 1433.410 2.400 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1468.270 -4.800 1468.830 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.210 -4.800 1486.770 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.690 -4.800 1504.250 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.050 -4.800 706.610 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1521.630 -4.800 1522.190 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.570 -4.800 1540.130 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1557.050 -4.800 1557.610 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1592.470 -4.800 1593.030 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.410 -4.800 1610.970 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.890 -4.800 1628.450 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1645.830 -4.800 1646.390 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1681.250 -4.800 1681.810 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 723.530 -4.800 724.090 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1716.670 -4.800 1717.230 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1734.610 -4.800 1735.170 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1752.090 -4.800 1752.650 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.030 -4.800 1770.590 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1805.450 -4.800 1806.010 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1822.930 -4.800 1823.490 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1840.870 -4.800 1841.430 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1858.350 -4.800 1858.910 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1876.290 -4.800 1876.850 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1894.230 -4.800 1894.790 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1929.650 -4.800 1930.210 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1982.550 -4.800 1983.110 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.490 -4.800 2001.050 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2017.970 -4.800 2018.530 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.950 -4.800 759.510 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2053.850 -4.800 2054.410 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.330 -4.800 2071.890 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2089.270 -4.800 2089.830 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2106.750 -4.800 2107.310 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.690 -4.800 2125.250 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2142.170 -4.800 2142.730 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2177.590 -4.800 2178.150 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 -4.800 2196.090 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2213.010 -4.800 2213.570 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 776.890 -4.800 777.450 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2230.950 -4.800 2231.510 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.890 -4.800 2249.450 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2266.370 -4.800 2266.930 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2301.790 -4.800 2302.350 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2319.730 -4.800 2320.290 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2337.210 -4.800 2337.770 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2355.150 -4.800 2355.710 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2390.570 -4.800 2391.130 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 794.370 -4.800 794.930 2.400 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.730 -4.800 641.290 2.400 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 2.400 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2431.970 -4.800 2432.530 2.400 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.450 -4.800 2450.010 2.400 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2467.390 -4.800 2467.950 2.400 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.330 -4.800 2485.890 2.400 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.810 -4.800 2503.370 2.400 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2520.750 -4.800 2521.310 2.400 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 2.400 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2556.170 -4.800 2556.730 2.400 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2573.650 -4.800 2574.210 2.400 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.290 -4.800 818.850 2.400 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2591.590 -4.800 2592.150 2.400 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.070 -4.800 2609.630 2.400 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2627.010 -4.800 2627.570 2.400 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2644.950 -4.800 2645.510 2.400 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 2.400 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2680.370 -4.800 2680.930 2.400 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2697.850 -4.800 2698.410 2.400 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2715.790 -4.800 2716.350 2.400 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2733.270 -4.800 2733.830 2.400 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2751.210 -4.800 2751.770 2.400 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.770 -4.800 836.330 2.400 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2768.690 -4.800 2769.250 2.400 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 2.400 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2804.110 -4.800 2804.670 2.400 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2822.050 -4.800 2822.610 2.400 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2839.990 -4.800 2840.550 2.400 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2857.470 -4.800 2858.030 2.400 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2875.410 -4.800 2875.970 2.400 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 853.710 -4.800 854.270 2.400 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 2.400 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 889.130 -4.800 889.690 2.400 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 2.400 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 924.550 -4.800 925.110 2.400 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.490 -4.800 943.050 2.400 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.970 -4.800 960.530 2.400 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 2.400 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 2.400 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1030.810 -4.800 1031.370 2.400 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1048.750 -4.800 1049.310 2.400 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1066.690 -4.800 1067.250 2.400 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1084.170 -4.800 1084.730 2.400 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1102.110 -4.800 1102.670 2.400 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 2.400 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1137.530 -4.800 1138.090 2.400 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.010 -4.800 1155.570 2.400 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.150 -4.800 676.710 2.400 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.950 -4.800 1173.510 2.400 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1190.430 -4.800 1190.990 2.400 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1208.370 -4.800 1208.930 2.400 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1225.850 -4.800 1226.410 2.400 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 2.400 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1261.730 -4.800 1262.290 2.400 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.210 -4.800 1279.770 2.400 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1297.150 -4.800 1297.710 2.400 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1314.630 -4.800 1315.190 2.400 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.570 -4.800 1333.130 2.400 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.090 -4.800 694.650 2.400 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1350.050 -4.800 1350.610 2.400 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 2.400 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1385.470 -4.800 1386.030 2.400 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.410 -4.800 1403.970 2.400 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1421.350 -4.800 1421.910 2.400 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1438.830 -4.800 1439.390 2.400 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.770 -4.800 1457.330 2.400 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1474.250 -4.800 1474.810 2.400 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 2.400 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1509.670 -4.800 1510.230 2.400 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 712.030 -4.800 712.590 2.400 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1527.610 -4.800 1528.170 2.400 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1545.090 -4.800 1545.650 2.400 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.030 -4.800 1563.590 2.400 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.970 -4.800 1581.530 2.400 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1598.450 -4.800 1599.010 2.400 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 2.400 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1633.870 -4.800 1634.430 2.400 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1651.810 -4.800 1652.370 2.400 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1669.290 -4.800 1669.850 2.400 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1687.230 -4.800 1687.790 2.400 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.510 -4.800 730.070 2.400 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 2.400 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1722.650 -4.800 1723.210 2.400 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.130 -4.800 1740.690 2.400 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.070 -4.800 1758.630 2.400 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.010 -4.800 1776.570 2.400 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.490 -4.800 1794.050 2.400 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1811.430 -4.800 1811.990 2.400 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 2.400 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1846.850 -4.800 1847.410 2.400 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.330 -4.800 1864.890 2.400 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 747.450 -4.800 748.010 2.400 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1882.270 -4.800 1882.830 2.400 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1935.630 -4.800 1936.190 2.400 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.530 -4.800 1989.090 2.400 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2023.950 -4.800 2024.510 2.400 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.890 -4.800 2042.450 2.400 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 764.930 -4.800 765.490 2.400 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2059.370 -4.800 2059.930 2.400 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 2.400 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2094.790 -4.800 2095.350 2.400 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2112.730 -4.800 2113.290 2.400 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2130.670 -4.800 2131.230 2.400 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2148.150 -4.800 2148.710 2.400 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2166.090 -4.800 2166.650 2.400 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 -4.800 2184.130 2.400 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 2.400 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.990 -4.800 2219.550 2.400 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 2.400 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2236.930 -4.800 2237.490 2.400 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2254.410 -4.800 2254.970 2.400 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2272.350 -4.800 2272.910 2.400 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2290.290 -4.800 2290.850 2.400 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2307.770 -4.800 2308.330 2.400 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 2.400 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2343.190 -4.800 2343.750 2.400 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.130 -4.800 2361.690 2.400 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.610 -4.800 2379.170 2.400 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.550 -4.800 2397.110 2.400 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.350 -4.800 800.910 2.400 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -10.030 -4.670 -6.930 3524.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 -4.670 2929.650 -1.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -10.030 3521.250 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2926.550 -4.670 2929.650 3524.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 23.970 -38.270 27.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 -38.270 91.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 407.145 91.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 683.145 91.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 959.145 91.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 1235.145 91.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 1511.145 91.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 1787.145 91.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 2063.145 91.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 2339.145 91.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 2615.145 91.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 2891.145 91.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 3167.145 91.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 88.470 3443.145 91.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 -38.270 156.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 407.145 156.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 683.145 156.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 959.145 156.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 1235.145 156.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 1511.145 156.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 1787.145 156.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 2063.145 156.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 2339.145 156.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 2615.145 156.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 2891.145 156.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 3167.145 156.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 152.970 3443.145 156.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 -38.270 220.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 407.145 220.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 683.145 220.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 959.145 220.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 1235.145 220.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 1511.145 220.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 1787.145 220.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 2063.145 220.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 2339.145 220.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 2615.145 220.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 2891.145 220.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 3167.145 220.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 217.470 3443.145 220.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 281.970 -38.270 285.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 -38.270 349.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 407.145 349.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 683.145 349.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 959.145 349.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 1235.145 349.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 1511.145 349.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 1787.145 349.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 2063.145 349.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 2339.145 349.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 2615.145 349.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 2891.145 349.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 3167.145 349.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 346.470 3443.145 349.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 -38.270 414.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 407.145 414.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 683.145 414.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 959.145 414.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 1235.145 414.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 1511.145 414.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 1787.145 414.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 2063.145 414.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 2339.145 414.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 2615.145 414.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 2891.145 414.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 3167.145 414.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 410.970 3443.145 414.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 -38.270 478.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 407.145 478.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 683.145 478.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 959.145 478.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 1235.145 478.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 1511.145 478.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 1787.145 478.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 2063.145 478.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 2339.145 478.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 2615.145 478.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 2891.145 478.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 3167.145 478.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 475.470 3443.145 478.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 539.970 -38.270 543.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 -38.270 607.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 407.145 607.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 683.145 607.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 959.145 607.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 1235.145 607.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 1511.145 607.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 1787.145 607.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 2063.145 607.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 2339.145 607.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 2615.145 607.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 2891.145 607.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 3167.145 607.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 604.470 3443.145 607.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 -38.270 672.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 407.145 672.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 683.145 672.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 959.145 672.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 1235.145 672.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 1511.145 672.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 1787.145 672.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 2063.145 672.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 2339.145 672.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 2615.145 672.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 2891.145 672.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 3167.145 672.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 668.970 3443.145 672.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 -38.270 736.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 407.145 736.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 683.145 736.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 959.145 736.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 1235.145 736.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 1511.145 736.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 1787.145 736.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 2063.145 736.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 2339.145 736.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 2615.145 736.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 2891.145 736.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 3167.145 736.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 733.470 3443.145 736.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 797.970 -38.270 801.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 -38.270 865.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 407.145 865.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 683.145 865.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 959.145 865.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 1235.145 865.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 1511.145 865.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 1787.145 865.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 2063.145 865.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 2339.145 865.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 2615.145 865.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 2891.145 865.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 3167.145 865.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 862.470 3443.145 865.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 -38.270 930.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 407.145 930.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 683.145 930.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 959.145 930.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 1235.145 930.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 1511.145 930.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 1787.145 930.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 2063.145 930.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 2339.145 930.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 2615.145 930.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 2891.145 930.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 3167.145 930.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 926.970 3443.145 930.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 -38.270 994.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 407.145 994.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 683.145 994.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 959.145 994.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 1235.145 994.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 1511.145 994.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 1787.145 994.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 2063.145 994.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 2339.145 994.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 2615.145 994.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 2891.145 994.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 3167.145 994.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 991.470 3443.145 994.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1055.970 -38.270 1059.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 -38.270 1123.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 407.145 1123.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 683.145 1123.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 959.145 1123.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 1235.145 1123.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 1511.145 1123.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 1787.145 1123.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 2063.145 1123.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 2339.145 1123.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 2615.145 1123.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 2891.145 1123.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 3167.145 1123.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1120.470 3443.145 1123.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 -38.270 1188.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 407.145 1188.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 683.145 1188.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 959.145 1188.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 1235.145 1188.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 1511.145 1188.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 1787.145 1188.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 2063.145 1188.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 2339.145 1188.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 2615.145 1188.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 2891.145 1188.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 3167.145 1188.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1184.970 3443.145 1188.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 -38.270 1252.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 407.145 1252.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 683.145 1252.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 959.145 1252.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 1235.145 1252.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 1511.145 1252.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 1787.145 1252.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 2063.145 1252.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 2339.145 1252.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 2615.145 1252.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 2891.145 1252.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 3167.145 1252.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.470 3443.145 1252.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1313.970 -38.270 1317.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 -38.270 1381.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 407.145 1381.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 683.145 1381.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 959.145 1381.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 1235.145 1381.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 1511.145 1381.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 1787.145 1381.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 2063.145 1381.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 2339.145 1381.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 2615.145 1381.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 2891.145 1381.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 3167.145 1381.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1378.470 3443.145 1381.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 -38.270 1446.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 407.145 1446.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 683.145 1446.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 959.145 1446.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 1235.145 1446.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 1511.145 1446.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 1787.145 1446.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 2063.145 1446.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 2339.145 1446.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 2615.145 1446.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 2891.145 1446.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 3167.145 1446.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1442.970 3443.145 1446.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 -38.270 1510.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 407.145 1510.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 683.145 1510.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 959.145 1510.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 1235.145 1510.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 1511.145 1510.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 1787.145 1510.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 2063.145 1510.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 2339.145 1510.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 2615.145 1510.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 2891.145 1510.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 3167.145 1510.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1507.470 3443.145 1510.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1571.970 -38.270 1575.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 -38.270 1639.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 407.145 1639.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 683.145 1639.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 959.145 1639.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 1235.145 1639.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 1511.145 1639.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 1787.145 1639.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 2063.145 1639.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 2339.145 1639.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 2615.145 1639.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 2891.145 1639.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 3167.145 1639.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1636.470 3443.145 1639.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 -38.270 1704.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 407.145 1704.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 683.145 1704.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 959.145 1704.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 1235.145 1704.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 1511.145 1704.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 1787.145 1704.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 2063.145 1704.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 2339.145 1704.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 2615.145 1704.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 2891.145 1704.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 3167.145 1704.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1700.970 3443.145 1704.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 -38.270 1768.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 407.145 1768.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 683.145 1768.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 959.145 1768.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 1235.145 1768.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 1511.145 1768.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 1787.145 1768.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 2063.145 1768.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 2339.145 1768.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 2615.145 1768.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 2891.145 1768.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 3167.145 1768.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1765.470 3443.145 1768.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1829.970 -38.270 1833.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 -38.270 1897.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 407.145 1897.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 683.145 1897.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 959.145 1897.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 1235.145 1897.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 1511.145 1897.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 1787.145 1897.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 2063.145 1897.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 2339.145 1897.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 2615.145 1897.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 2891.145 1897.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 3167.145 1897.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1894.470 3443.145 1897.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 -38.270 1962.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 407.145 1962.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 683.145 1962.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 959.145 1962.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 1235.145 1962.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 1511.145 1962.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 1787.145 1962.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 2063.145 1962.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 2339.145 1962.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 2615.145 1962.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 2891.145 1962.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 3167.145 1962.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1958.970 3443.145 1962.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 -38.270 2026.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 407.145 2026.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 683.145 2026.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 959.145 2026.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 1235.145 2026.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 1511.145 2026.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 1787.145 2026.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 2063.145 2026.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 2339.145 2026.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 2615.145 2026.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 2891.145 2026.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 3167.145 2026.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2023.470 3443.145 2026.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2087.970 -38.270 2091.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 -38.270 2155.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 407.145 2155.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 683.145 2155.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 959.145 2155.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 1235.145 2155.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 1511.145 2155.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 1787.145 2155.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 2063.145 2155.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 2339.145 2155.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 2615.145 2155.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 2891.145 2155.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 3167.145 2155.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2152.470 3443.145 2155.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 -38.270 2220.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 407.145 2220.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 683.145 2220.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 959.145 2220.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 1235.145 2220.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 1511.145 2220.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 1787.145 2220.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 2063.145 2220.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 2339.145 2220.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 2615.145 2220.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 2891.145 2220.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 3167.145 2220.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2216.970 3443.145 2220.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 -38.270 2284.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 407.145 2284.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 683.145 2284.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 959.145 2284.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 1235.145 2284.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 1511.145 2284.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 1787.145 2284.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 2063.145 2284.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 2339.145 2284.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 2615.145 2284.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 2891.145 2284.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 3167.145 2284.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2281.470 3443.145 2284.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2345.970 -38.270 2349.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 -38.270 2413.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 407.145 2413.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 683.145 2413.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 959.145 2413.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 1235.145 2413.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 1511.145 2413.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 1787.145 2413.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 2063.145 2413.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 2339.145 2413.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 2615.145 2413.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 2891.145 2413.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 3167.145 2413.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2410.470 3443.145 2413.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 -38.270 2478.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 407.145 2478.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 683.145 2478.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 959.145 2478.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 1235.145 2478.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 1511.145 2478.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 1787.145 2478.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 2063.145 2478.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 2339.145 2478.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 2615.145 2478.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 2891.145 2478.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 3167.145 2478.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2474.970 3443.145 2478.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 -38.270 2542.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 407.145 2542.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 683.145 2542.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 959.145 2542.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 1235.145 2542.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 1511.145 2542.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 1787.145 2542.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 2063.145 2542.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 2339.145 2542.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 2615.145 2542.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 2891.145 2542.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 3167.145 2542.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2539.470 3443.145 2542.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2603.970 -38.270 2607.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 -38.270 2671.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 407.145 2671.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 683.145 2671.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 959.145 2671.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 1235.145 2671.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 1511.145 2671.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 1787.145 2671.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 2063.145 2671.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 2339.145 2671.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 2615.145 2671.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 2891.145 2671.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 3167.145 2671.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2668.470 3443.145 2671.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 -38.270 2736.070 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 407.145 2736.070 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 683.145 2736.070 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 959.145 2736.070 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 1235.145 2736.070 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 1511.145 2736.070 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 1787.145 2736.070 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 2063.145 2736.070 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 2339.145 2736.070 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 2615.145 2736.070 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 2891.145 2736.070 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 3167.145 2736.070 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2732.970 3443.145 2736.070 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 -38.270 2800.570 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 407.145 2800.570 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 683.145 2800.570 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 959.145 2800.570 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 1235.145 2800.570 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 1511.145 2800.570 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 1787.145 2800.570 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 2063.145 2800.570 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 2339.145 2800.570 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 2615.145 2800.570 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 2891.145 2800.570 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 3167.145 2800.570 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2797.470 3443.145 2800.570 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2861.970 -38.270 2865.070 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 49.330 2963.250 52.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 83.830 2963.250 86.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 118.330 2963.250 121.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 152.830 2963.250 155.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 187.330 2963.250 190.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 221.830 2963.250 224.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 256.330 2963.250 259.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 290.830 2963.250 293.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 325.330 2963.250 328.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 359.830 2963.250 362.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 394.330 2963.250 397.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 428.830 2963.250 431.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 463.330 2963.250 466.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 497.830 2963.250 500.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 532.330 2963.250 535.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 566.830 2963.250 569.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 601.330 2963.250 604.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 635.830 2963.250 638.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 670.330 2963.250 673.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 704.830 2963.250 707.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 739.330 2963.250 742.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 773.830 2963.250 776.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 808.330 2963.250 811.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 842.830 2963.250 845.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 877.330 2963.250 880.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 911.830 2963.250 914.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 946.330 2963.250 949.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 980.830 2963.250 983.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1015.330 2963.250 1018.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1049.830 2963.250 1052.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1084.330 2963.250 1087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1118.830 2963.250 1121.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1153.330 2963.250 1156.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1187.830 2963.250 1190.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1222.330 2963.250 1225.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1256.830 2963.250 1259.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1291.330 2963.250 1294.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1325.830 2963.250 1328.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1360.330 2963.250 1363.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1394.830 2963.250 1397.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1429.330 2963.250 1432.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1463.830 2963.250 1466.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1498.330 2963.250 1501.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1532.830 2963.250 1535.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1567.330 2963.250 1570.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1601.830 2963.250 1604.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1636.330 2963.250 1639.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1670.830 2963.250 1673.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1705.330 2963.250 1708.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1739.830 2963.250 1742.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1774.330 2963.250 1777.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1808.830 2963.250 1811.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1843.330 2963.250 1846.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1877.830 2963.250 1880.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1912.330 2963.250 1915.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1946.830 2963.250 1949.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1981.330 2963.250 1984.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2015.830 2963.250 2018.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2050.330 2963.250 2053.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2084.830 2963.250 2087.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2119.330 2963.250 2122.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2153.830 2963.250 2156.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2188.330 2963.250 2191.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2222.830 2963.250 2225.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2257.330 2963.250 2260.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2291.830 2963.250 2294.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2326.330 2963.250 2329.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2360.830 2963.250 2363.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2395.330 2963.250 2398.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2429.830 2963.250 2432.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2464.330 2963.250 2467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2498.830 2963.250 2501.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2533.330 2963.250 2536.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2567.830 2963.250 2570.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2602.330 2963.250 2605.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2636.830 2963.250 2639.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2671.330 2963.250 2674.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2705.830 2963.250 2708.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2740.330 2963.250 2743.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2774.830 2963.250 2777.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2809.330 2963.250 2812.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2843.830 2963.250 2846.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2878.330 2963.250 2881.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2912.830 2963.250 2915.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2947.330 2963.250 2950.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2981.830 2963.250 2984.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3016.330 2963.250 3019.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3050.830 2963.250 3053.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3085.330 2963.250 3088.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3119.830 2963.250 3122.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3154.330 2963.250 3157.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3188.830 2963.250 3191.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3223.330 2963.250 3226.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3257.830 2963.250 3260.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3292.330 2963.250 3295.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3326.830 2963.250 3329.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3361.330 2963.250 3364.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3395.830 2963.250 3398.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3430.330 2963.250 3433.430 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3464.830 2963.250 3467.930 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3499.330 2963.250 3502.430 ;
    END
  END vccd1
  PIN vccd2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -19.630 -14.270 -16.530 3533.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 -14.270 2939.250 -11.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -19.630 3530.850 2939.250 3533.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2936.150 -14.270 2939.250 3533.950 ;
    END
  END vccd2
  PIN vdda1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -29.230 -23.870 -26.130 3543.550 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 -23.870 2948.850 -20.770 ;
    END
    PORT
      LAYER met5 ;
        RECT -29.230 3540.450 2948.850 3543.550 ;
    END
    PORT
      LAYER met4 ;
        RECT 2945.750 -23.870 2948.850 3543.550 ;
    END
  END vdda1
  PIN vdda2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT -38.830 -33.470 -35.730 3553.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 -33.470 2958.450 -30.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -38.830 3550.050 2958.450 3553.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2955.350 -33.470 2958.450 3553.150 ;
    END
  END vdda2
  PIN vssa1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -34.030 -28.670 -30.930 3548.350 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 -28.670 2953.650 -25.570 ;
    END
    PORT
      LAYER met5 ;
        RECT -34.030 3545.250 2953.650 3548.350 ;
    END
    PORT
      LAYER met4 ;
        RECT 2950.550 -28.670 2953.650 3548.350 ;
    END
  END vssa1
  PIN vssa2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -43.630 -38.270 -40.530 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 -38.270 2963.250 -35.170 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3554.850 2963.250 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2960.150 -38.270 2963.250 3557.950 ;
    END
  END vssa2
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -14.830 -9.470 -11.730 3529.150 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 -9.470 2934.450 -6.370 ;
    END
    PORT
      LAYER met5 ;
        RECT -14.830 3526.050 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 2931.350 -9.470 2934.450 3529.150 ;
    END
    PORT
      LAYER met4 ;
        RECT 56.220 -38.270 59.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 -38.270 123.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 407.145 123.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 683.145 123.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 959.145 123.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 1235.145 123.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 1511.145 123.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 1787.145 123.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 2063.145 123.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 2339.145 123.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 2615.145 123.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 2891.145 123.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 3167.145 123.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 120.720 3443.145 123.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 -38.270 188.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 407.145 188.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 683.145 188.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 959.145 188.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 1235.145 188.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 1511.145 188.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 1787.145 188.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 2063.145 188.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 2339.145 188.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 2615.145 188.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 2891.145 188.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 3167.145 188.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 185.220 3443.145 188.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 -38.270 252.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 407.145 252.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 683.145 252.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 959.145 252.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 1235.145 252.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 1511.145 252.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 1787.145 252.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 2063.145 252.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 2339.145 252.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 2615.145 252.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 2891.145 252.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 3167.145 252.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.720 3443.145 252.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 314.220 -38.270 317.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 -38.270 381.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 407.145 381.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 683.145 381.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 959.145 381.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 1235.145 381.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 1511.145 381.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 1787.145 381.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 2063.145 381.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 2339.145 381.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 2615.145 381.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 2891.145 381.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 3167.145 381.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 378.720 3443.145 381.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 -38.270 446.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 407.145 446.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 683.145 446.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 959.145 446.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 1235.145 446.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 1511.145 446.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 1787.145 446.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 2063.145 446.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 2339.145 446.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 2615.145 446.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 2891.145 446.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 3167.145 446.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 443.220 3443.145 446.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 -38.270 510.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 407.145 510.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 683.145 510.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 959.145 510.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 1235.145 510.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 1511.145 510.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 1787.145 510.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 2063.145 510.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 2339.145 510.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 2615.145 510.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 2891.145 510.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 3167.145 510.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 507.720 3443.145 510.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 572.220 -38.270 575.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 -38.270 639.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 407.145 639.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 683.145 639.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 959.145 639.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 1235.145 639.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 1511.145 639.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 1787.145 639.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 2063.145 639.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 2339.145 639.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 2615.145 639.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 2891.145 639.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 3167.145 639.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 636.720 3443.145 639.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 -38.270 704.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 407.145 704.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 683.145 704.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 959.145 704.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 1235.145 704.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 1511.145 704.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 1787.145 704.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 2063.145 704.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 2339.145 704.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 2615.145 704.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 2891.145 704.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 3167.145 704.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 701.220 3443.145 704.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 -38.270 768.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 407.145 768.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 683.145 768.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 959.145 768.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 1235.145 768.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 1511.145 768.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 1787.145 768.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 2063.145 768.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 2339.145 768.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 2615.145 768.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 2891.145 768.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 3167.145 768.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 765.720 3443.145 768.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 830.220 -38.270 833.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 -38.270 897.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 407.145 897.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 683.145 897.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 959.145 897.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 1235.145 897.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 1511.145 897.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 1787.145 897.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 2063.145 897.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 2339.145 897.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 2615.145 897.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 2891.145 897.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 3167.145 897.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 894.720 3443.145 897.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 -38.270 962.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 407.145 962.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 683.145 962.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 959.145 962.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 1235.145 962.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 1511.145 962.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 1787.145 962.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 2063.145 962.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 2339.145 962.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 2615.145 962.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 2891.145 962.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 3167.145 962.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 959.220 3443.145 962.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 -38.270 1026.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 407.145 1026.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 683.145 1026.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 959.145 1026.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 1235.145 1026.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 1511.145 1026.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 1787.145 1026.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 2063.145 1026.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 2339.145 1026.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 2615.145 1026.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 2891.145 1026.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 3167.145 1026.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1023.720 3443.145 1026.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.220 -38.270 1091.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 -38.270 1155.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 407.145 1155.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 683.145 1155.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 959.145 1155.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 1235.145 1155.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 1511.145 1155.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 1787.145 1155.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 2063.145 1155.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 2339.145 1155.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 2615.145 1155.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 2891.145 1155.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 3167.145 1155.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1152.720 3443.145 1155.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 -38.270 1220.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 407.145 1220.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 683.145 1220.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 959.145 1220.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 1235.145 1220.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 1511.145 1220.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 1787.145 1220.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 2063.145 1220.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 2339.145 1220.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 2615.145 1220.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 2891.145 1220.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 3167.145 1220.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1217.220 3443.145 1220.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 -38.270 1284.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 407.145 1284.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 683.145 1284.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 959.145 1284.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 1235.145 1284.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 1511.145 1284.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 1787.145 1284.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 2063.145 1284.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 2339.145 1284.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 2615.145 1284.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 2891.145 1284.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 3167.145 1284.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1281.720 3443.145 1284.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1346.220 -38.270 1349.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 -38.270 1413.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 407.145 1413.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 683.145 1413.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 959.145 1413.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 1235.145 1413.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 1511.145 1413.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 1787.145 1413.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 2063.145 1413.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 2339.145 1413.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 2615.145 1413.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 2891.145 1413.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 3167.145 1413.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1410.720 3443.145 1413.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 -38.270 1478.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 407.145 1478.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 683.145 1478.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 959.145 1478.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 1235.145 1478.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 1511.145 1478.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 1787.145 1478.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 2063.145 1478.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 2339.145 1478.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 2615.145 1478.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 2891.145 1478.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 3167.145 1478.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1475.220 3443.145 1478.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 -38.270 1542.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 407.145 1542.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 683.145 1542.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 959.145 1542.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 1235.145 1542.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 1511.145 1542.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 1787.145 1542.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 2063.145 1542.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 2339.145 1542.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 2615.145 1542.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 2891.145 1542.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 3167.145 1542.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1539.720 3443.145 1542.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1604.220 -38.270 1607.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 -38.270 1671.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 407.145 1671.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 683.145 1671.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 959.145 1671.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 1235.145 1671.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 1511.145 1671.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 1787.145 1671.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 2063.145 1671.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 2339.145 1671.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 2615.145 1671.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 2891.145 1671.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 3167.145 1671.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1668.720 3443.145 1671.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 -38.270 1736.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 407.145 1736.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 683.145 1736.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 959.145 1736.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 1235.145 1736.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 1511.145 1736.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 1787.145 1736.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 2063.145 1736.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 2339.145 1736.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 2615.145 1736.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 2891.145 1736.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 3167.145 1736.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1733.220 3443.145 1736.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 -38.270 1800.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 407.145 1800.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 683.145 1800.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 959.145 1800.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 1235.145 1800.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 1511.145 1800.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 1787.145 1800.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 2063.145 1800.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 2339.145 1800.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 2615.145 1800.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 2891.145 1800.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 3167.145 1800.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1797.720 3443.145 1800.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1862.220 -38.270 1865.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 -38.270 1929.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 407.145 1929.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 683.145 1929.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 959.145 1929.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 1235.145 1929.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 1511.145 1929.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 1787.145 1929.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 2063.145 1929.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 2339.145 1929.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 2615.145 1929.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 2891.145 1929.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 3167.145 1929.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1926.720 3443.145 1929.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 -38.270 1994.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 407.145 1994.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 683.145 1994.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 959.145 1994.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 1235.145 1994.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 1511.145 1994.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 1787.145 1994.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 2063.145 1994.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 2339.145 1994.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 2615.145 1994.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 2891.145 1994.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 3167.145 1994.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1991.220 3443.145 1994.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 -38.270 2058.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 407.145 2058.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 683.145 2058.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 959.145 2058.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 1235.145 2058.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 1511.145 2058.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 1787.145 2058.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 2063.145 2058.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 2339.145 2058.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 2615.145 2058.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 2891.145 2058.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 3167.145 2058.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2055.720 3443.145 2058.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2120.220 -38.270 2123.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 -38.270 2187.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 407.145 2187.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 683.145 2187.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 959.145 2187.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 1235.145 2187.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 1511.145 2187.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 1787.145 2187.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 2063.145 2187.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 2339.145 2187.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 2615.145 2187.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 2891.145 2187.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 3167.145 2187.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2184.720 3443.145 2187.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 -38.270 2252.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 407.145 2252.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 683.145 2252.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 959.145 2252.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 1235.145 2252.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 1511.145 2252.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 1787.145 2252.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 2063.145 2252.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 2339.145 2252.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 2615.145 2252.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 2891.145 2252.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 3167.145 2252.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2249.220 3443.145 2252.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 -38.270 2316.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 407.145 2316.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 683.145 2316.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 959.145 2316.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 1235.145 2316.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 1511.145 2316.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 1787.145 2316.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 2063.145 2316.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 2339.145 2316.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 2615.145 2316.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 2891.145 2316.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 3167.145 2316.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2313.720 3443.145 2316.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2378.220 -38.270 2381.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 -38.270 2445.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 407.145 2445.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 683.145 2445.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 959.145 2445.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 1235.145 2445.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 1511.145 2445.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 1787.145 2445.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 2063.145 2445.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 2339.145 2445.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 2615.145 2445.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 2891.145 2445.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 3167.145 2445.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2442.720 3443.145 2445.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 -38.270 2510.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 407.145 2510.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 683.145 2510.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 959.145 2510.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 1235.145 2510.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 1511.145 2510.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 1787.145 2510.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 2063.145 2510.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 2339.145 2510.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 2615.145 2510.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 2891.145 2510.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 3167.145 2510.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2507.220 3443.145 2510.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 -38.270 2574.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 407.145 2574.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 683.145 2574.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 959.145 2574.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 1235.145 2574.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 1511.145 2574.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 1787.145 2574.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 2063.145 2574.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 2339.145 2574.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 2615.145 2574.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 2891.145 2574.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 3167.145 2574.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2571.720 3443.145 2574.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2636.220 -38.270 2639.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 -38.270 2703.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 407.145 2703.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 683.145 2703.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 959.145 2703.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 1235.145 2703.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 1511.145 2703.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 1787.145 2703.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 2063.145 2703.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 2339.145 2703.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 2615.145 2703.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 2891.145 2703.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 3167.145 2703.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2700.720 3443.145 2703.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 -38.270 2768.320 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 407.145 2768.320 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 683.145 2768.320 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 959.145 2768.320 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 1235.145 2768.320 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 1511.145 2768.320 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 1787.145 2768.320 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 2063.145 2768.320 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 2339.145 2768.320 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 2615.145 2768.320 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 2891.145 2768.320 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 3167.145 2768.320 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2765.220 3443.145 2768.320 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 -38.270 2832.820 190.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 407.145 2832.820 466.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 683.145 2832.820 742.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 959.145 2832.820 1018.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 1235.145 2832.820 1294.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 1511.145 2832.820 1570.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 1787.145 2832.820 1846.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 2063.145 2832.820 2122.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 2339.145 2832.820 2398.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 2615.145 2832.820 2674.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 2891.145 2832.820 2950.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 3167.145 2832.820 3226.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2829.720 3443.145 2832.820 3557.950 ;
    END
    PORT
      LAYER met4 ;
        RECT 2894.220 -38.270 2897.320 3557.950 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 66.580 2963.250 69.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 101.080 2963.250 104.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 135.580 2963.250 138.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 170.080 2963.250 173.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 204.580 2963.250 207.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 239.080 2963.250 242.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 273.580 2963.250 276.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 308.080 2963.250 311.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 342.580 2963.250 345.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 377.080 2963.250 380.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 411.580 2963.250 414.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 446.080 2963.250 449.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 480.580 2963.250 483.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 515.080 2963.250 518.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 549.580 2963.250 552.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 584.080 2963.250 587.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 618.580 2963.250 621.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 653.080 2963.250 656.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 687.580 2963.250 690.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 722.080 2963.250 725.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 756.580 2963.250 759.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 791.080 2963.250 794.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 825.580 2963.250 828.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 860.080 2963.250 863.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 894.580 2963.250 897.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 929.080 2963.250 932.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 963.580 2963.250 966.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 998.080 2963.250 1001.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1032.580 2963.250 1035.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1067.080 2963.250 1070.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1101.580 2963.250 1104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1136.080 2963.250 1139.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1170.580 2963.250 1173.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1205.080 2963.250 1208.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1239.580 2963.250 1242.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1274.080 2963.250 1277.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1308.580 2963.250 1311.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1343.080 2963.250 1346.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1377.580 2963.250 1380.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1412.080 2963.250 1415.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1446.580 2963.250 1449.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1481.080 2963.250 1484.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1515.580 2963.250 1518.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1550.080 2963.250 1553.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1584.580 2963.250 1587.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1619.080 2963.250 1622.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1653.580 2963.250 1656.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1688.080 2963.250 1691.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1722.580 2963.250 1725.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1757.080 2963.250 1760.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1791.580 2963.250 1794.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1826.080 2963.250 1829.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1860.580 2963.250 1863.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1895.080 2963.250 1898.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1929.580 2963.250 1932.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1964.080 2963.250 1967.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 1998.580 2963.250 2001.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2033.080 2963.250 2036.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2067.580 2963.250 2070.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2102.080 2963.250 2105.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2136.580 2963.250 2139.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2171.080 2963.250 2174.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2205.580 2963.250 2208.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2240.080 2963.250 2243.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2274.580 2963.250 2277.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2309.080 2963.250 2312.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2343.580 2963.250 2346.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2378.080 2963.250 2381.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2412.580 2963.250 2415.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2447.080 2963.250 2450.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2481.580 2963.250 2484.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2516.080 2963.250 2519.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2550.580 2963.250 2553.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2585.080 2963.250 2588.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2619.580 2963.250 2622.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2654.080 2963.250 2657.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2688.580 2963.250 2691.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2723.080 2963.250 2726.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2757.580 2963.250 2760.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2792.080 2963.250 2795.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2826.580 2963.250 2829.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2861.080 2963.250 2864.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2895.580 2963.250 2898.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2930.080 2963.250 2933.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2964.580 2963.250 2967.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 2999.080 2963.250 3002.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3033.580 2963.250 3036.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3068.080 2963.250 3071.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3102.580 2963.250 3105.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3137.080 2963.250 3140.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3171.580 2963.250 3174.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3206.080 2963.250 3209.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3240.580 2963.250 3243.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3275.080 2963.250 3278.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3309.580 2963.250 3312.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3344.080 2963.250 3347.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3378.580 2963.250 3381.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3413.080 2963.250 3416.180 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3447.580 2963.250 3450.680 ;
    END
    PORT
      LAYER met5 ;
        RECT -43.630 3482.080 2963.250 3485.180 ;
    END
  END vssd1
  PIN vssd2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT -24.430 -19.070 -21.330 3538.750 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 -19.070 2944.050 -15.970 ;
    END
    PORT
      LAYER met5 ;
        RECT -24.430 3535.650 2944.050 3538.750 ;
    END
    PORT
      LAYER met4 ;
        RECT 2940.950 -19.070 2944.050 3538.750 ;
    END
  END vssd2
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 256.630 -4.800 257.190 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.570 -4.800 275.130 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.050 -4.800 292.610 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.990 -4.800 310.550 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 345.410 -4.800 345.970 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 362.890 -4.800 363.450 2.400 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.830 -4.800 381.390 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 398.310 -4.800 398.870 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.590 -4.800 62.150 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 416.250 -4.800 416.810 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.190 -4.800 434.750 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 469.610 -4.800 470.170 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.090 -4.800 487.650 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.030 -4.800 505.590 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.510 -4.800 523.070 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 540.450 -4.800 541.010 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.930 -4.800 558.490 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.050 -4.800 85.610 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.810 -4.800 594.370 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.290 -4.800 611.850 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.970 -4.800 109.530 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.430 -4.800 132.990 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.370 -4.800 150.930 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.850 -4.800 168.410 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 185.790 -4.800 186.350 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.210 -4.800 221.770 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 20.190 -4.800 20.750 2.400 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 43.650 -4.800 44.210 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.610 -4.800 263.170 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.090 -4.800 280.650 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.030 -4.800 298.590 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.970 -4.800 316.530 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.450 -4.800 334.010 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.390 -4.800 351.950 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.810 -4.800 387.370 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.290 -4.800 404.850 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.570 -4.800 68.130 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 422.230 -4.800 422.790 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 439.710 -4.800 440.270 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.650 -4.800 458.210 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.590 -4.800 476.150 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 511.010 -4.800 511.570 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.490 -4.800 529.050 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.430 -4.800 546.990 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.910 -4.800 564.470 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.850 -4.800 582.410 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 91.030 -4.800 91.590 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 599.330 -4.800 599.890 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.410 -4.800 138.970 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.830 -4.800 174.390 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.770 -4.800 192.330 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.250 -4.800 209.810 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 227.190 -4.800 227.750 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.630 -4.800 50.190 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.650 -4.800 251.210 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 268.590 -4.800 269.150 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.010 -4.800 304.570 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.490 -4.800 322.050 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 339.430 -4.800 339.990 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.370 -4.800 357.930 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.850 -4.800 375.410 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.790 -4.800 393.350 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 2.400 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.550 -4.800 74.110 2.400 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.210 -4.800 428.770 2.400 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 445.690 -4.800 446.250 2.400 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 463.630 -4.800 464.190 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 481.110 -4.800 481.670 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.050 -4.800 499.610 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 516.530 -4.800 517.090 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.410 -4.800 552.970 2.400 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.890 -4.800 570.450 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 587.830 -4.800 588.390 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.010 -4.800 97.570 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 605.310 -4.800 605.870 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 623.250 -4.800 623.810 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.930 -4.800 121.490 2.400 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.390 -4.800 144.950 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 2.400 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.810 -4.800 180.370 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.230 -4.800 215.790 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.170 -4.800 233.730 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.610 -4.800 56.170 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.530 -4.800 80.090 2.400 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.990 -4.800 103.550 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 -4.800 127.010 2.400 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.150 -4.800 32.710 2.400 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2914.100 3508.885 ;
      LAYER met1 ;
        RECT 4.210 3.780 2917.250 3512.840 ;
      LAYER met2 ;
        RECT 0.550 3517.320 40.150 3518.050 ;
        RECT 41.270 3517.320 121.110 3518.050 ;
        RECT 122.230 3517.320 202.070 3518.050 ;
        RECT 203.190 3517.320 283.490 3518.050 ;
        RECT 284.610 3517.320 364.450 3518.050 ;
        RECT 365.570 3517.320 445.410 3518.050 ;
        RECT 446.530 3517.320 526.830 3518.050 ;
        RECT 527.950 3517.320 607.790 3518.050 ;
        RECT 608.910 3517.320 688.750 3518.050 ;
        RECT 689.870 3517.320 770.170 3518.050 ;
        RECT 771.290 3517.320 851.130 3518.050 ;
        RECT 852.250 3517.320 932.090 3518.050 ;
        RECT 933.210 3517.320 1013.510 3518.050 ;
        RECT 1014.630 3517.320 1094.470 3518.050 ;
        RECT 1095.590 3517.320 1175.430 3518.050 ;
        RECT 1176.550 3517.320 1256.850 3518.050 ;
        RECT 1257.970 3517.320 1337.810 3518.050 ;
        RECT 1338.930 3517.320 1418.770 3518.050 ;
        RECT 1419.890 3517.320 1500.190 3518.050 ;
        RECT 1501.310 3517.320 1581.150 3518.050 ;
        RECT 1582.270 3517.320 1662.110 3518.050 ;
        RECT 1663.230 3517.320 1743.530 3518.050 ;
        RECT 1744.650 3517.320 1824.490 3518.050 ;
        RECT 1825.610 3517.320 1905.450 3518.050 ;
        RECT 1906.570 3517.320 1986.870 3518.050 ;
        RECT 1987.990 3517.320 2067.830 3518.050 ;
        RECT 2068.950 3517.320 2148.790 3518.050 ;
        RECT 2149.910 3517.320 2230.210 3518.050 ;
        RECT 2231.330 3517.320 2311.170 3518.050 ;
        RECT 2312.290 3517.320 2392.130 3518.050 ;
        RECT 2393.250 3517.320 2473.550 3518.050 ;
        RECT 2474.670 3517.320 2554.510 3518.050 ;
        RECT 2555.630 3517.320 2635.470 3518.050 ;
        RECT 2636.590 3517.320 2716.890 3518.050 ;
        RECT 2718.010 3517.320 2797.850 3518.050 ;
        RECT 2798.970 3517.320 2878.810 3518.050 ;
        RECT 2879.930 3517.320 2917.220 3518.050 ;
        RECT 0.550 2.680 2917.220 3517.320 ;
        RECT 0.550 0.155 2.430 2.680 ;
        RECT 3.550 0.155 7.950 2.680 ;
        RECT 9.070 0.155 13.930 2.680 ;
        RECT 15.050 0.155 19.910 2.680 ;
        RECT 21.030 0.155 25.890 2.680 ;
        RECT 27.010 0.155 31.870 2.680 ;
        RECT 32.990 0.155 37.850 2.680 ;
        RECT 38.970 0.155 43.370 2.680 ;
        RECT 44.490 0.155 49.350 2.680 ;
        RECT 50.470 0.155 55.330 2.680 ;
        RECT 56.450 0.155 61.310 2.680 ;
        RECT 62.430 0.155 67.290 2.680 ;
        RECT 68.410 0.155 73.270 2.680 ;
        RECT 74.390 0.155 79.250 2.680 ;
        RECT 80.370 0.155 84.770 2.680 ;
        RECT 85.890 0.155 90.750 2.680 ;
        RECT 91.870 0.155 96.730 2.680 ;
        RECT 97.850 0.155 102.710 2.680 ;
        RECT 103.830 0.155 108.690 2.680 ;
        RECT 109.810 0.155 114.670 2.680 ;
        RECT 115.790 0.155 120.650 2.680 ;
        RECT 121.770 0.155 126.170 2.680 ;
        RECT 127.290 0.155 132.150 2.680 ;
        RECT 133.270 0.155 138.130 2.680 ;
        RECT 139.250 0.155 144.110 2.680 ;
        RECT 145.230 0.155 150.090 2.680 ;
        RECT 151.210 0.155 156.070 2.680 ;
        RECT 157.190 0.155 161.590 2.680 ;
        RECT 162.710 0.155 167.570 2.680 ;
        RECT 168.690 0.155 173.550 2.680 ;
        RECT 174.670 0.155 179.530 2.680 ;
        RECT 180.650 0.155 185.510 2.680 ;
        RECT 186.630 0.155 191.490 2.680 ;
        RECT 192.610 0.155 197.470 2.680 ;
        RECT 198.590 0.155 202.990 2.680 ;
        RECT 204.110 0.155 208.970 2.680 ;
        RECT 210.090 0.155 214.950 2.680 ;
        RECT 216.070 0.155 220.930 2.680 ;
        RECT 222.050 0.155 226.910 2.680 ;
        RECT 228.030 0.155 232.890 2.680 ;
        RECT 234.010 0.155 238.870 2.680 ;
        RECT 239.990 0.155 244.390 2.680 ;
        RECT 245.510 0.155 250.370 2.680 ;
        RECT 251.490 0.155 256.350 2.680 ;
        RECT 257.470 0.155 262.330 2.680 ;
        RECT 263.450 0.155 268.310 2.680 ;
        RECT 269.430 0.155 274.290 2.680 ;
        RECT 275.410 0.155 279.810 2.680 ;
        RECT 280.930 0.155 285.790 2.680 ;
        RECT 286.910 0.155 291.770 2.680 ;
        RECT 292.890 0.155 297.750 2.680 ;
        RECT 298.870 0.155 303.730 2.680 ;
        RECT 304.850 0.155 309.710 2.680 ;
        RECT 310.830 0.155 315.690 2.680 ;
        RECT 316.810 0.155 321.210 2.680 ;
        RECT 322.330 0.155 327.190 2.680 ;
        RECT 328.310 0.155 333.170 2.680 ;
        RECT 334.290 0.155 339.150 2.680 ;
        RECT 340.270 0.155 345.130 2.680 ;
        RECT 346.250 0.155 351.110 2.680 ;
        RECT 352.230 0.155 357.090 2.680 ;
        RECT 358.210 0.155 362.610 2.680 ;
        RECT 363.730 0.155 368.590 2.680 ;
        RECT 369.710 0.155 374.570 2.680 ;
        RECT 375.690 0.155 380.550 2.680 ;
        RECT 381.670 0.155 386.530 2.680 ;
        RECT 387.650 0.155 392.510 2.680 ;
        RECT 393.630 0.155 398.030 2.680 ;
        RECT 399.150 0.155 404.010 2.680 ;
        RECT 405.130 0.155 409.990 2.680 ;
        RECT 411.110 0.155 415.970 2.680 ;
        RECT 417.090 0.155 421.950 2.680 ;
        RECT 423.070 0.155 427.930 2.680 ;
        RECT 429.050 0.155 433.910 2.680 ;
        RECT 435.030 0.155 439.430 2.680 ;
        RECT 440.550 0.155 445.410 2.680 ;
        RECT 446.530 0.155 451.390 2.680 ;
        RECT 452.510 0.155 457.370 2.680 ;
        RECT 458.490 0.155 463.350 2.680 ;
        RECT 464.470 0.155 469.330 2.680 ;
        RECT 470.450 0.155 475.310 2.680 ;
        RECT 476.430 0.155 480.830 2.680 ;
        RECT 481.950 0.155 486.810 2.680 ;
        RECT 487.930 0.155 492.790 2.680 ;
        RECT 493.910 0.155 498.770 2.680 ;
        RECT 499.890 0.155 504.750 2.680 ;
        RECT 505.870 0.155 510.730 2.680 ;
        RECT 511.850 0.155 516.250 2.680 ;
        RECT 517.370 0.155 522.230 2.680 ;
        RECT 523.350 0.155 528.210 2.680 ;
        RECT 529.330 0.155 534.190 2.680 ;
        RECT 535.310 0.155 540.170 2.680 ;
        RECT 541.290 0.155 546.150 2.680 ;
        RECT 547.270 0.155 552.130 2.680 ;
        RECT 553.250 0.155 557.650 2.680 ;
        RECT 558.770 0.155 563.630 2.680 ;
        RECT 564.750 0.155 569.610 2.680 ;
        RECT 570.730 0.155 575.590 2.680 ;
        RECT 576.710 0.155 581.570 2.680 ;
        RECT 582.690 0.155 587.550 2.680 ;
        RECT 588.670 0.155 593.530 2.680 ;
        RECT 594.650 0.155 599.050 2.680 ;
        RECT 600.170 0.155 605.030 2.680 ;
        RECT 606.150 0.155 611.010 2.680 ;
        RECT 612.130 0.155 616.990 2.680 ;
        RECT 618.110 0.155 622.970 2.680 ;
        RECT 624.090 0.155 628.950 2.680 ;
        RECT 630.070 0.155 634.470 2.680 ;
        RECT 635.590 0.155 640.450 2.680 ;
        RECT 641.570 0.155 646.430 2.680 ;
        RECT 647.550 0.155 652.410 2.680 ;
        RECT 653.530 0.155 658.390 2.680 ;
        RECT 659.510 0.155 664.370 2.680 ;
        RECT 665.490 0.155 670.350 2.680 ;
        RECT 671.470 0.155 675.870 2.680 ;
        RECT 676.990 0.155 681.850 2.680 ;
        RECT 682.970 0.155 687.830 2.680 ;
        RECT 688.950 0.155 693.810 2.680 ;
        RECT 694.930 0.155 699.790 2.680 ;
        RECT 700.910 0.155 705.770 2.680 ;
        RECT 706.890 0.155 711.750 2.680 ;
        RECT 712.870 0.155 717.270 2.680 ;
        RECT 718.390 0.155 723.250 2.680 ;
        RECT 724.370 0.155 729.230 2.680 ;
        RECT 730.350 0.155 735.210 2.680 ;
        RECT 736.330 0.155 741.190 2.680 ;
        RECT 742.310 0.155 747.170 2.680 ;
        RECT 748.290 0.155 752.690 2.680 ;
        RECT 753.810 0.155 758.670 2.680 ;
        RECT 759.790 0.155 764.650 2.680 ;
        RECT 765.770 0.155 770.630 2.680 ;
        RECT 771.750 0.155 776.610 2.680 ;
        RECT 777.730 0.155 782.590 2.680 ;
        RECT 783.710 0.155 788.570 2.680 ;
        RECT 789.690 0.155 794.090 2.680 ;
        RECT 795.210 0.155 800.070 2.680 ;
        RECT 801.190 0.155 806.050 2.680 ;
        RECT 807.170 0.155 812.030 2.680 ;
        RECT 813.150 0.155 818.010 2.680 ;
        RECT 819.130 0.155 823.990 2.680 ;
        RECT 825.110 0.155 829.970 2.680 ;
        RECT 831.090 0.155 835.490 2.680 ;
        RECT 836.610 0.155 841.470 2.680 ;
        RECT 842.590 0.155 847.450 2.680 ;
        RECT 848.570 0.155 853.430 2.680 ;
        RECT 854.550 0.155 859.410 2.680 ;
        RECT 860.530 0.155 865.390 2.680 ;
        RECT 866.510 0.155 870.910 2.680 ;
        RECT 872.030 0.155 876.890 2.680 ;
        RECT 878.010 0.155 882.870 2.680 ;
        RECT 883.990 0.155 888.850 2.680 ;
        RECT 889.970 0.155 894.830 2.680 ;
        RECT 895.950 0.155 900.810 2.680 ;
        RECT 901.930 0.155 906.790 2.680 ;
        RECT 907.910 0.155 912.310 2.680 ;
        RECT 913.430 0.155 918.290 2.680 ;
        RECT 919.410 0.155 924.270 2.680 ;
        RECT 925.390 0.155 930.250 2.680 ;
        RECT 931.370 0.155 936.230 2.680 ;
        RECT 937.350 0.155 942.210 2.680 ;
        RECT 943.330 0.155 948.190 2.680 ;
        RECT 949.310 0.155 953.710 2.680 ;
        RECT 954.830 0.155 959.690 2.680 ;
        RECT 960.810 0.155 965.670 2.680 ;
        RECT 966.790 0.155 971.650 2.680 ;
        RECT 972.770 0.155 977.630 2.680 ;
        RECT 978.750 0.155 983.610 2.680 ;
        RECT 984.730 0.155 989.130 2.680 ;
        RECT 990.250 0.155 995.110 2.680 ;
        RECT 996.230 0.155 1001.090 2.680 ;
        RECT 1002.210 0.155 1007.070 2.680 ;
        RECT 1008.190 0.155 1013.050 2.680 ;
        RECT 1014.170 0.155 1019.030 2.680 ;
        RECT 1020.150 0.155 1025.010 2.680 ;
        RECT 1026.130 0.155 1030.530 2.680 ;
        RECT 1031.650 0.155 1036.510 2.680 ;
        RECT 1037.630 0.155 1042.490 2.680 ;
        RECT 1043.610 0.155 1048.470 2.680 ;
        RECT 1049.590 0.155 1054.450 2.680 ;
        RECT 1055.570 0.155 1060.430 2.680 ;
        RECT 1061.550 0.155 1066.410 2.680 ;
        RECT 1067.530 0.155 1071.930 2.680 ;
        RECT 1073.050 0.155 1077.910 2.680 ;
        RECT 1079.030 0.155 1083.890 2.680 ;
        RECT 1085.010 0.155 1089.870 2.680 ;
        RECT 1090.990 0.155 1095.850 2.680 ;
        RECT 1096.970 0.155 1101.830 2.680 ;
        RECT 1102.950 0.155 1107.350 2.680 ;
        RECT 1108.470 0.155 1113.330 2.680 ;
        RECT 1114.450 0.155 1119.310 2.680 ;
        RECT 1120.430 0.155 1125.290 2.680 ;
        RECT 1126.410 0.155 1131.270 2.680 ;
        RECT 1132.390 0.155 1137.250 2.680 ;
        RECT 1138.370 0.155 1143.230 2.680 ;
        RECT 1144.350 0.155 1148.750 2.680 ;
        RECT 1149.870 0.155 1154.730 2.680 ;
        RECT 1155.850 0.155 1160.710 2.680 ;
        RECT 1161.830 0.155 1166.690 2.680 ;
        RECT 1167.810 0.155 1172.670 2.680 ;
        RECT 1173.790 0.155 1178.650 2.680 ;
        RECT 1179.770 0.155 1184.630 2.680 ;
        RECT 1185.750 0.155 1190.150 2.680 ;
        RECT 1191.270 0.155 1196.130 2.680 ;
        RECT 1197.250 0.155 1202.110 2.680 ;
        RECT 1203.230 0.155 1208.090 2.680 ;
        RECT 1209.210 0.155 1214.070 2.680 ;
        RECT 1215.190 0.155 1220.050 2.680 ;
        RECT 1221.170 0.155 1225.570 2.680 ;
        RECT 1226.690 0.155 1231.550 2.680 ;
        RECT 1232.670 0.155 1237.530 2.680 ;
        RECT 1238.650 0.155 1243.510 2.680 ;
        RECT 1244.630 0.155 1249.490 2.680 ;
        RECT 1250.610 0.155 1255.470 2.680 ;
        RECT 1256.590 0.155 1261.450 2.680 ;
        RECT 1262.570 0.155 1266.970 2.680 ;
        RECT 1268.090 0.155 1272.950 2.680 ;
        RECT 1274.070 0.155 1278.930 2.680 ;
        RECT 1280.050 0.155 1284.910 2.680 ;
        RECT 1286.030 0.155 1290.890 2.680 ;
        RECT 1292.010 0.155 1296.870 2.680 ;
        RECT 1297.990 0.155 1302.850 2.680 ;
        RECT 1303.970 0.155 1308.370 2.680 ;
        RECT 1309.490 0.155 1314.350 2.680 ;
        RECT 1315.470 0.155 1320.330 2.680 ;
        RECT 1321.450 0.155 1326.310 2.680 ;
        RECT 1327.430 0.155 1332.290 2.680 ;
        RECT 1333.410 0.155 1338.270 2.680 ;
        RECT 1339.390 0.155 1343.790 2.680 ;
        RECT 1344.910 0.155 1349.770 2.680 ;
        RECT 1350.890 0.155 1355.750 2.680 ;
        RECT 1356.870 0.155 1361.730 2.680 ;
        RECT 1362.850 0.155 1367.710 2.680 ;
        RECT 1368.830 0.155 1373.690 2.680 ;
        RECT 1374.810 0.155 1379.670 2.680 ;
        RECT 1380.790 0.155 1385.190 2.680 ;
        RECT 1386.310 0.155 1391.170 2.680 ;
        RECT 1392.290 0.155 1397.150 2.680 ;
        RECT 1398.270 0.155 1403.130 2.680 ;
        RECT 1404.250 0.155 1409.110 2.680 ;
        RECT 1410.230 0.155 1415.090 2.680 ;
        RECT 1416.210 0.155 1421.070 2.680 ;
        RECT 1422.190 0.155 1426.590 2.680 ;
        RECT 1427.710 0.155 1432.570 2.680 ;
        RECT 1433.690 0.155 1438.550 2.680 ;
        RECT 1439.670 0.155 1444.530 2.680 ;
        RECT 1445.650 0.155 1450.510 2.680 ;
        RECT 1451.630 0.155 1456.490 2.680 ;
        RECT 1457.610 0.155 1462.470 2.680 ;
        RECT 1463.590 0.155 1467.990 2.680 ;
        RECT 1469.110 0.155 1473.970 2.680 ;
        RECT 1475.090 0.155 1479.950 2.680 ;
        RECT 1481.070 0.155 1485.930 2.680 ;
        RECT 1487.050 0.155 1491.910 2.680 ;
        RECT 1493.030 0.155 1497.890 2.680 ;
        RECT 1499.010 0.155 1503.410 2.680 ;
        RECT 1504.530 0.155 1509.390 2.680 ;
        RECT 1510.510 0.155 1515.370 2.680 ;
        RECT 1516.490 0.155 1521.350 2.680 ;
        RECT 1522.470 0.155 1527.330 2.680 ;
        RECT 1528.450 0.155 1533.310 2.680 ;
        RECT 1534.430 0.155 1539.290 2.680 ;
        RECT 1540.410 0.155 1544.810 2.680 ;
        RECT 1545.930 0.155 1550.790 2.680 ;
        RECT 1551.910 0.155 1556.770 2.680 ;
        RECT 1557.890 0.155 1562.750 2.680 ;
        RECT 1563.870 0.155 1568.730 2.680 ;
        RECT 1569.850 0.155 1574.710 2.680 ;
        RECT 1575.830 0.155 1580.690 2.680 ;
        RECT 1581.810 0.155 1586.210 2.680 ;
        RECT 1587.330 0.155 1592.190 2.680 ;
        RECT 1593.310 0.155 1598.170 2.680 ;
        RECT 1599.290 0.155 1604.150 2.680 ;
        RECT 1605.270 0.155 1610.130 2.680 ;
        RECT 1611.250 0.155 1616.110 2.680 ;
        RECT 1617.230 0.155 1621.630 2.680 ;
        RECT 1622.750 0.155 1627.610 2.680 ;
        RECT 1628.730 0.155 1633.590 2.680 ;
        RECT 1634.710 0.155 1639.570 2.680 ;
        RECT 1640.690 0.155 1645.550 2.680 ;
        RECT 1646.670 0.155 1651.530 2.680 ;
        RECT 1652.650 0.155 1657.510 2.680 ;
        RECT 1658.630 0.155 1663.030 2.680 ;
        RECT 1664.150 0.155 1669.010 2.680 ;
        RECT 1670.130 0.155 1674.990 2.680 ;
        RECT 1676.110 0.155 1680.970 2.680 ;
        RECT 1682.090 0.155 1686.950 2.680 ;
        RECT 1688.070 0.155 1692.930 2.680 ;
        RECT 1694.050 0.155 1698.910 2.680 ;
        RECT 1700.030 0.155 1704.430 2.680 ;
        RECT 1705.550 0.155 1710.410 2.680 ;
        RECT 1711.530 0.155 1716.390 2.680 ;
        RECT 1717.510 0.155 1722.370 2.680 ;
        RECT 1723.490 0.155 1728.350 2.680 ;
        RECT 1729.470 0.155 1734.330 2.680 ;
        RECT 1735.450 0.155 1739.850 2.680 ;
        RECT 1740.970 0.155 1745.830 2.680 ;
        RECT 1746.950 0.155 1751.810 2.680 ;
        RECT 1752.930 0.155 1757.790 2.680 ;
        RECT 1758.910 0.155 1763.770 2.680 ;
        RECT 1764.890 0.155 1769.750 2.680 ;
        RECT 1770.870 0.155 1775.730 2.680 ;
        RECT 1776.850 0.155 1781.250 2.680 ;
        RECT 1782.370 0.155 1787.230 2.680 ;
        RECT 1788.350 0.155 1793.210 2.680 ;
        RECT 1794.330 0.155 1799.190 2.680 ;
        RECT 1800.310 0.155 1805.170 2.680 ;
        RECT 1806.290 0.155 1811.150 2.680 ;
        RECT 1812.270 0.155 1817.130 2.680 ;
        RECT 1818.250 0.155 1822.650 2.680 ;
        RECT 1823.770 0.155 1828.630 2.680 ;
        RECT 1829.750 0.155 1834.610 2.680 ;
        RECT 1835.730 0.155 1840.590 2.680 ;
        RECT 1841.710 0.155 1846.570 2.680 ;
        RECT 1847.690 0.155 1852.550 2.680 ;
        RECT 1853.670 0.155 1858.070 2.680 ;
        RECT 1859.190 0.155 1864.050 2.680 ;
        RECT 1865.170 0.155 1870.030 2.680 ;
        RECT 1871.150 0.155 1876.010 2.680 ;
        RECT 1877.130 0.155 1881.990 2.680 ;
        RECT 1883.110 0.155 1887.970 2.680 ;
        RECT 1889.090 0.155 1893.950 2.680 ;
        RECT 1895.070 0.155 1899.470 2.680 ;
        RECT 1900.590 0.155 1905.450 2.680 ;
        RECT 1906.570 0.155 1911.430 2.680 ;
        RECT 1912.550 0.155 1917.410 2.680 ;
        RECT 1918.530 0.155 1923.390 2.680 ;
        RECT 1924.510 0.155 1929.370 2.680 ;
        RECT 1930.490 0.155 1935.350 2.680 ;
        RECT 1936.470 0.155 1940.870 2.680 ;
        RECT 1941.990 0.155 1946.850 2.680 ;
        RECT 1947.970 0.155 1952.830 2.680 ;
        RECT 1953.950 0.155 1958.810 2.680 ;
        RECT 1959.930 0.155 1964.790 2.680 ;
        RECT 1965.910 0.155 1970.770 2.680 ;
        RECT 1971.890 0.155 1976.290 2.680 ;
        RECT 1977.410 0.155 1982.270 2.680 ;
        RECT 1983.390 0.155 1988.250 2.680 ;
        RECT 1989.370 0.155 1994.230 2.680 ;
        RECT 1995.350 0.155 2000.210 2.680 ;
        RECT 2001.330 0.155 2006.190 2.680 ;
        RECT 2007.310 0.155 2012.170 2.680 ;
        RECT 2013.290 0.155 2017.690 2.680 ;
        RECT 2018.810 0.155 2023.670 2.680 ;
        RECT 2024.790 0.155 2029.650 2.680 ;
        RECT 2030.770 0.155 2035.630 2.680 ;
        RECT 2036.750 0.155 2041.610 2.680 ;
        RECT 2042.730 0.155 2047.590 2.680 ;
        RECT 2048.710 0.155 2053.570 2.680 ;
        RECT 2054.690 0.155 2059.090 2.680 ;
        RECT 2060.210 0.155 2065.070 2.680 ;
        RECT 2066.190 0.155 2071.050 2.680 ;
        RECT 2072.170 0.155 2077.030 2.680 ;
        RECT 2078.150 0.155 2083.010 2.680 ;
        RECT 2084.130 0.155 2088.990 2.680 ;
        RECT 2090.110 0.155 2094.510 2.680 ;
        RECT 2095.630 0.155 2100.490 2.680 ;
        RECT 2101.610 0.155 2106.470 2.680 ;
        RECT 2107.590 0.155 2112.450 2.680 ;
        RECT 2113.570 0.155 2118.430 2.680 ;
        RECT 2119.550 0.155 2124.410 2.680 ;
        RECT 2125.530 0.155 2130.390 2.680 ;
        RECT 2131.510 0.155 2135.910 2.680 ;
        RECT 2137.030 0.155 2141.890 2.680 ;
        RECT 2143.010 0.155 2147.870 2.680 ;
        RECT 2148.990 0.155 2153.850 2.680 ;
        RECT 2154.970 0.155 2159.830 2.680 ;
        RECT 2160.950 0.155 2165.810 2.680 ;
        RECT 2166.930 0.155 2171.790 2.680 ;
        RECT 2172.910 0.155 2177.310 2.680 ;
        RECT 2178.430 0.155 2183.290 2.680 ;
        RECT 2184.410 0.155 2189.270 2.680 ;
        RECT 2190.390 0.155 2195.250 2.680 ;
        RECT 2196.370 0.155 2201.230 2.680 ;
        RECT 2202.350 0.155 2207.210 2.680 ;
        RECT 2208.330 0.155 2212.730 2.680 ;
        RECT 2213.850 0.155 2218.710 2.680 ;
        RECT 2219.830 0.155 2224.690 2.680 ;
        RECT 2225.810 0.155 2230.670 2.680 ;
        RECT 2231.790 0.155 2236.650 2.680 ;
        RECT 2237.770 0.155 2242.630 2.680 ;
        RECT 2243.750 0.155 2248.610 2.680 ;
        RECT 2249.730 0.155 2254.130 2.680 ;
        RECT 2255.250 0.155 2260.110 2.680 ;
        RECT 2261.230 0.155 2266.090 2.680 ;
        RECT 2267.210 0.155 2272.070 2.680 ;
        RECT 2273.190 0.155 2278.050 2.680 ;
        RECT 2279.170 0.155 2284.030 2.680 ;
        RECT 2285.150 0.155 2290.010 2.680 ;
        RECT 2291.130 0.155 2295.530 2.680 ;
        RECT 2296.650 0.155 2301.510 2.680 ;
        RECT 2302.630 0.155 2307.490 2.680 ;
        RECT 2308.610 0.155 2313.470 2.680 ;
        RECT 2314.590 0.155 2319.450 2.680 ;
        RECT 2320.570 0.155 2325.430 2.680 ;
        RECT 2326.550 0.155 2330.950 2.680 ;
        RECT 2332.070 0.155 2336.930 2.680 ;
        RECT 2338.050 0.155 2342.910 2.680 ;
        RECT 2344.030 0.155 2348.890 2.680 ;
        RECT 2350.010 0.155 2354.870 2.680 ;
        RECT 2355.990 0.155 2360.850 2.680 ;
        RECT 2361.970 0.155 2366.830 2.680 ;
        RECT 2367.950 0.155 2372.350 2.680 ;
        RECT 2373.470 0.155 2378.330 2.680 ;
        RECT 2379.450 0.155 2384.310 2.680 ;
        RECT 2385.430 0.155 2390.290 2.680 ;
        RECT 2391.410 0.155 2396.270 2.680 ;
        RECT 2397.390 0.155 2402.250 2.680 ;
        RECT 2403.370 0.155 2408.230 2.680 ;
        RECT 2409.350 0.155 2413.750 2.680 ;
        RECT 2414.870 0.155 2419.730 2.680 ;
        RECT 2420.850 0.155 2425.710 2.680 ;
        RECT 2426.830 0.155 2431.690 2.680 ;
        RECT 2432.810 0.155 2437.670 2.680 ;
        RECT 2438.790 0.155 2443.650 2.680 ;
        RECT 2444.770 0.155 2449.170 2.680 ;
        RECT 2450.290 0.155 2455.150 2.680 ;
        RECT 2456.270 0.155 2461.130 2.680 ;
        RECT 2462.250 0.155 2467.110 2.680 ;
        RECT 2468.230 0.155 2473.090 2.680 ;
        RECT 2474.210 0.155 2479.070 2.680 ;
        RECT 2480.190 0.155 2485.050 2.680 ;
        RECT 2486.170 0.155 2490.570 2.680 ;
        RECT 2491.690 0.155 2496.550 2.680 ;
        RECT 2497.670 0.155 2502.530 2.680 ;
        RECT 2503.650 0.155 2508.510 2.680 ;
        RECT 2509.630 0.155 2514.490 2.680 ;
        RECT 2515.610 0.155 2520.470 2.680 ;
        RECT 2521.590 0.155 2526.450 2.680 ;
        RECT 2527.570 0.155 2531.970 2.680 ;
        RECT 2533.090 0.155 2537.950 2.680 ;
        RECT 2539.070 0.155 2543.930 2.680 ;
        RECT 2545.050 0.155 2549.910 2.680 ;
        RECT 2551.030 0.155 2555.890 2.680 ;
        RECT 2557.010 0.155 2561.870 2.680 ;
        RECT 2562.990 0.155 2567.390 2.680 ;
        RECT 2568.510 0.155 2573.370 2.680 ;
        RECT 2574.490 0.155 2579.350 2.680 ;
        RECT 2580.470 0.155 2585.330 2.680 ;
        RECT 2586.450 0.155 2591.310 2.680 ;
        RECT 2592.430 0.155 2597.290 2.680 ;
        RECT 2598.410 0.155 2603.270 2.680 ;
        RECT 2604.390 0.155 2608.790 2.680 ;
        RECT 2609.910 0.155 2614.770 2.680 ;
        RECT 2615.890 0.155 2620.750 2.680 ;
        RECT 2621.870 0.155 2626.730 2.680 ;
        RECT 2627.850 0.155 2632.710 2.680 ;
        RECT 2633.830 0.155 2638.690 2.680 ;
        RECT 2639.810 0.155 2644.670 2.680 ;
        RECT 2645.790 0.155 2650.190 2.680 ;
        RECT 2651.310 0.155 2656.170 2.680 ;
        RECT 2657.290 0.155 2662.150 2.680 ;
        RECT 2663.270 0.155 2668.130 2.680 ;
        RECT 2669.250 0.155 2674.110 2.680 ;
        RECT 2675.230 0.155 2680.090 2.680 ;
        RECT 2681.210 0.155 2685.610 2.680 ;
        RECT 2686.730 0.155 2691.590 2.680 ;
        RECT 2692.710 0.155 2697.570 2.680 ;
        RECT 2698.690 0.155 2703.550 2.680 ;
        RECT 2704.670 0.155 2709.530 2.680 ;
        RECT 2710.650 0.155 2715.510 2.680 ;
        RECT 2716.630 0.155 2721.490 2.680 ;
        RECT 2722.610 0.155 2727.010 2.680 ;
        RECT 2728.130 0.155 2732.990 2.680 ;
        RECT 2734.110 0.155 2738.970 2.680 ;
        RECT 2740.090 0.155 2744.950 2.680 ;
        RECT 2746.070 0.155 2750.930 2.680 ;
        RECT 2752.050 0.155 2756.910 2.680 ;
        RECT 2758.030 0.155 2762.890 2.680 ;
        RECT 2764.010 0.155 2768.410 2.680 ;
        RECT 2769.530 0.155 2774.390 2.680 ;
        RECT 2775.510 0.155 2780.370 2.680 ;
        RECT 2781.490 0.155 2786.350 2.680 ;
        RECT 2787.470 0.155 2792.330 2.680 ;
        RECT 2793.450 0.155 2798.310 2.680 ;
        RECT 2799.430 0.155 2803.830 2.680 ;
        RECT 2804.950 0.155 2809.810 2.680 ;
        RECT 2810.930 0.155 2815.790 2.680 ;
        RECT 2816.910 0.155 2821.770 2.680 ;
        RECT 2822.890 0.155 2827.750 2.680 ;
        RECT 2828.870 0.155 2833.730 2.680 ;
        RECT 2834.850 0.155 2839.710 2.680 ;
        RECT 2840.830 0.155 2845.230 2.680 ;
        RECT 2846.350 0.155 2851.210 2.680 ;
        RECT 2852.330 0.155 2857.190 2.680 ;
        RECT 2858.310 0.155 2863.170 2.680 ;
        RECT 2864.290 0.155 2869.150 2.680 ;
        RECT 2870.270 0.155 2875.130 2.680 ;
        RECT 2876.250 0.155 2881.110 2.680 ;
        RECT 2882.230 0.155 2886.630 2.680 ;
        RECT 2887.750 0.155 2892.610 2.680 ;
        RECT 2893.730 0.155 2898.590 2.680 ;
        RECT 2899.710 0.155 2904.570 2.680 ;
        RECT 2905.690 0.155 2910.550 2.680 ;
        RECT 2911.670 0.155 2916.530 2.680 ;
      LAYER met3 ;
        RECT 0.525 3487.700 2917.600 3512.700 ;
        RECT 2.800 3487.020 2917.600 3487.700 ;
        RECT 2.800 3485.700 2917.200 3487.020 ;
        RECT 0.525 3485.020 2917.200 3485.700 ;
        RECT 0.525 3422.420 2917.600 3485.020 ;
        RECT 2.800 3420.420 2917.600 3422.420 ;
        RECT 0.525 3420.380 2917.600 3420.420 ;
        RECT 0.525 3418.380 2917.200 3420.380 ;
        RECT 0.525 3357.140 2917.600 3418.380 ;
        RECT 2.800 3355.140 2917.600 3357.140 ;
        RECT 0.525 3354.420 2917.600 3355.140 ;
        RECT 0.525 3352.420 2917.200 3354.420 ;
        RECT 0.525 3291.860 2917.600 3352.420 ;
        RECT 2.800 3289.860 2917.600 3291.860 ;
        RECT 0.525 3287.780 2917.600 3289.860 ;
        RECT 0.525 3285.780 2917.200 3287.780 ;
        RECT 0.525 3226.580 2917.600 3285.780 ;
        RECT 2.800 3224.580 2917.600 3226.580 ;
        RECT 0.525 3221.140 2917.600 3224.580 ;
        RECT 0.525 3219.140 2917.200 3221.140 ;
        RECT 0.525 3161.300 2917.600 3219.140 ;
        RECT 2.800 3159.300 2917.600 3161.300 ;
        RECT 0.525 3155.180 2917.600 3159.300 ;
        RECT 0.525 3153.180 2917.200 3155.180 ;
        RECT 0.525 3096.700 2917.600 3153.180 ;
        RECT 2.800 3094.700 2917.600 3096.700 ;
        RECT 0.525 3088.540 2917.600 3094.700 ;
        RECT 0.525 3086.540 2917.200 3088.540 ;
        RECT 0.525 3031.420 2917.600 3086.540 ;
        RECT 2.800 3029.420 2917.600 3031.420 ;
        RECT 0.525 3021.900 2917.600 3029.420 ;
        RECT 0.525 3019.900 2917.200 3021.900 ;
        RECT 0.525 2966.140 2917.600 3019.900 ;
        RECT 2.800 2964.140 2917.600 2966.140 ;
        RECT 0.525 2955.940 2917.600 2964.140 ;
        RECT 0.525 2953.940 2917.200 2955.940 ;
        RECT 0.525 2900.860 2917.600 2953.940 ;
        RECT 2.800 2898.860 2917.600 2900.860 ;
        RECT 0.525 2889.300 2917.600 2898.860 ;
        RECT 0.525 2887.300 2917.200 2889.300 ;
        RECT 0.525 2835.580 2917.600 2887.300 ;
        RECT 2.800 2833.580 2917.600 2835.580 ;
        RECT 0.525 2822.660 2917.600 2833.580 ;
        RECT 0.525 2820.660 2917.200 2822.660 ;
        RECT 0.525 2770.300 2917.600 2820.660 ;
        RECT 2.800 2768.300 2917.600 2770.300 ;
        RECT 0.525 2756.700 2917.600 2768.300 ;
        RECT 0.525 2754.700 2917.200 2756.700 ;
        RECT 0.525 2705.020 2917.600 2754.700 ;
        RECT 2.800 2703.020 2917.600 2705.020 ;
        RECT 0.525 2690.060 2917.600 2703.020 ;
        RECT 0.525 2688.060 2917.200 2690.060 ;
        RECT 0.525 2640.420 2917.600 2688.060 ;
        RECT 2.800 2638.420 2917.600 2640.420 ;
        RECT 0.525 2623.420 2917.600 2638.420 ;
        RECT 0.525 2621.420 2917.200 2623.420 ;
        RECT 0.525 2575.140 2917.600 2621.420 ;
        RECT 2.800 2573.140 2917.600 2575.140 ;
        RECT 0.525 2557.460 2917.600 2573.140 ;
        RECT 0.525 2555.460 2917.200 2557.460 ;
        RECT 0.525 2509.860 2917.600 2555.460 ;
        RECT 2.800 2507.860 2917.600 2509.860 ;
        RECT 0.525 2490.820 2917.600 2507.860 ;
        RECT 0.525 2488.820 2917.200 2490.820 ;
        RECT 0.525 2444.580 2917.600 2488.820 ;
        RECT 2.800 2442.580 2917.600 2444.580 ;
        RECT 0.525 2424.180 2917.600 2442.580 ;
        RECT 0.525 2422.180 2917.200 2424.180 ;
        RECT 0.525 2379.300 2917.600 2422.180 ;
        RECT 2.800 2377.300 2917.600 2379.300 ;
        RECT 0.525 2358.220 2917.600 2377.300 ;
        RECT 0.525 2356.220 2917.200 2358.220 ;
        RECT 0.525 2314.020 2917.600 2356.220 ;
        RECT 2.800 2312.020 2917.600 2314.020 ;
        RECT 0.525 2291.580 2917.600 2312.020 ;
        RECT 0.525 2289.580 2917.200 2291.580 ;
        RECT 0.525 2248.740 2917.600 2289.580 ;
        RECT 2.800 2246.740 2917.600 2248.740 ;
        RECT 0.525 2224.940 2917.600 2246.740 ;
        RECT 0.525 2222.940 2917.200 2224.940 ;
        RECT 0.525 2184.140 2917.600 2222.940 ;
        RECT 2.800 2182.140 2917.600 2184.140 ;
        RECT 0.525 2158.980 2917.600 2182.140 ;
        RECT 0.525 2156.980 2917.200 2158.980 ;
        RECT 0.525 2118.860 2917.600 2156.980 ;
        RECT 2.800 2116.860 2917.600 2118.860 ;
        RECT 0.525 2092.340 2917.600 2116.860 ;
        RECT 0.525 2090.340 2917.200 2092.340 ;
        RECT 0.525 2053.580 2917.600 2090.340 ;
        RECT 2.800 2051.580 2917.600 2053.580 ;
        RECT 0.525 2025.700 2917.600 2051.580 ;
        RECT 0.525 2023.700 2917.200 2025.700 ;
        RECT 0.525 1988.300 2917.600 2023.700 ;
        RECT 2.800 1986.300 2917.600 1988.300 ;
        RECT 0.525 1959.740 2917.600 1986.300 ;
        RECT 0.525 1957.740 2917.200 1959.740 ;
        RECT 0.525 1923.020 2917.600 1957.740 ;
        RECT 2.800 1921.020 2917.600 1923.020 ;
        RECT 0.525 1893.100 2917.600 1921.020 ;
        RECT 0.525 1891.100 2917.200 1893.100 ;
        RECT 0.525 1857.740 2917.600 1891.100 ;
        RECT 2.800 1855.740 2917.600 1857.740 ;
        RECT 0.525 1826.460 2917.600 1855.740 ;
        RECT 0.525 1824.460 2917.200 1826.460 ;
        RECT 0.525 1793.140 2917.600 1824.460 ;
        RECT 2.800 1791.140 2917.600 1793.140 ;
        RECT 0.525 1760.500 2917.600 1791.140 ;
        RECT 0.525 1758.500 2917.200 1760.500 ;
        RECT 0.525 1727.860 2917.600 1758.500 ;
        RECT 2.800 1725.860 2917.600 1727.860 ;
        RECT 0.525 1693.860 2917.600 1725.860 ;
        RECT 0.525 1691.860 2917.200 1693.860 ;
        RECT 0.525 1662.580 2917.600 1691.860 ;
        RECT 2.800 1660.580 2917.600 1662.580 ;
        RECT 0.525 1627.220 2917.600 1660.580 ;
        RECT 0.525 1625.220 2917.200 1627.220 ;
        RECT 0.525 1597.300 2917.600 1625.220 ;
        RECT 2.800 1595.300 2917.600 1597.300 ;
        RECT 0.525 1561.260 2917.600 1595.300 ;
        RECT 0.525 1559.260 2917.200 1561.260 ;
        RECT 0.525 1532.020 2917.600 1559.260 ;
        RECT 2.800 1530.020 2917.600 1532.020 ;
        RECT 0.525 1494.620 2917.600 1530.020 ;
        RECT 0.525 1492.620 2917.200 1494.620 ;
        RECT 0.525 1466.740 2917.600 1492.620 ;
        RECT 2.800 1464.740 2917.600 1466.740 ;
        RECT 0.525 1427.980 2917.600 1464.740 ;
        RECT 0.525 1425.980 2917.200 1427.980 ;
        RECT 0.525 1401.460 2917.600 1425.980 ;
        RECT 2.800 1399.460 2917.600 1401.460 ;
        RECT 0.525 1362.020 2917.600 1399.460 ;
        RECT 0.525 1360.020 2917.200 1362.020 ;
        RECT 0.525 1336.860 2917.600 1360.020 ;
        RECT 2.800 1334.860 2917.600 1336.860 ;
        RECT 0.525 1295.380 2917.600 1334.860 ;
        RECT 0.525 1293.380 2917.200 1295.380 ;
        RECT 0.525 1271.580 2917.600 1293.380 ;
        RECT 2.800 1269.580 2917.600 1271.580 ;
        RECT 0.525 1228.740 2917.600 1269.580 ;
        RECT 0.525 1226.740 2917.200 1228.740 ;
        RECT 0.525 1206.300 2917.600 1226.740 ;
        RECT 2.800 1204.300 2917.600 1206.300 ;
        RECT 0.525 1162.780 2917.600 1204.300 ;
        RECT 0.525 1160.780 2917.200 1162.780 ;
        RECT 0.525 1141.020 2917.600 1160.780 ;
        RECT 2.800 1139.020 2917.600 1141.020 ;
        RECT 0.525 1096.140 2917.600 1139.020 ;
        RECT 0.525 1094.140 2917.200 1096.140 ;
        RECT 0.525 1075.740 2917.600 1094.140 ;
        RECT 2.800 1073.740 2917.600 1075.740 ;
        RECT 0.525 1029.500 2917.600 1073.740 ;
        RECT 0.525 1027.500 2917.200 1029.500 ;
        RECT 0.525 1010.460 2917.600 1027.500 ;
        RECT 2.800 1008.460 2917.600 1010.460 ;
        RECT 0.525 963.540 2917.600 1008.460 ;
        RECT 0.525 961.540 2917.200 963.540 ;
        RECT 0.525 945.180 2917.600 961.540 ;
        RECT 2.800 943.180 2917.600 945.180 ;
        RECT 0.525 896.900 2917.600 943.180 ;
        RECT 0.525 894.900 2917.200 896.900 ;
        RECT 0.525 880.580 2917.600 894.900 ;
        RECT 2.800 878.580 2917.600 880.580 ;
        RECT 0.525 830.260 2917.600 878.580 ;
        RECT 0.525 828.260 2917.200 830.260 ;
        RECT 0.525 815.300 2917.600 828.260 ;
        RECT 2.800 813.300 2917.600 815.300 ;
        RECT 0.525 764.300 2917.600 813.300 ;
        RECT 0.525 762.300 2917.200 764.300 ;
        RECT 0.525 750.020 2917.600 762.300 ;
        RECT 2.800 748.020 2917.600 750.020 ;
        RECT 0.525 697.660 2917.600 748.020 ;
        RECT 0.525 695.660 2917.200 697.660 ;
        RECT 0.525 684.740 2917.600 695.660 ;
        RECT 2.800 682.740 2917.600 684.740 ;
        RECT 0.525 631.020 2917.600 682.740 ;
        RECT 0.525 629.020 2917.200 631.020 ;
        RECT 0.525 619.460 2917.600 629.020 ;
        RECT 2.800 617.460 2917.600 619.460 ;
        RECT 0.525 565.060 2917.600 617.460 ;
        RECT 0.525 563.060 2917.200 565.060 ;
        RECT 0.525 554.180 2917.600 563.060 ;
        RECT 2.800 552.180 2917.600 554.180 ;
        RECT 0.525 498.420 2917.600 552.180 ;
        RECT 0.525 496.420 2917.200 498.420 ;
        RECT 0.525 488.900 2917.600 496.420 ;
        RECT 2.800 486.900 2917.600 488.900 ;
        RECT 0.525 431.780 2917.600 486.900 ;
        RECT 0.525 429.780 2917.200 431.780 ;
        RECT 0.525 424.300 2917.600 429.780 ;
        RECT 2.800 422.300 2917.600 424.300 ;
        RECT 0.525 365.820 2917.600 422.300 ;
        RECT 0.525 363.820 2917.200 365.820 ;
        RECT 0.525 359.020 2917.600 363.820 ;
        RECT 2.800 357.020 2917.600 359.020 ;
        RECT 0.525 299.180 2917.600 357.020 ;
        RECT 0.525 297.180 2917.200 299.180 ;
        RECT 0.525 293.740 2917.600 297.180 ;
        RECT 2.800 291.740 2917.600 293.740 ;
        RECT 0.525 232.540 2917.600 291.740 ;
        RECT 0.525 230.540 2917.200 232.540 ;
        RECT 0.525 228.460 2917.600 230.540 ;
        RECT 2.800 226.460 2917.600 228.460 ;
        RECT 0.525 166.580 2917.600 226.460 ;
        RECT 0.525 164.580 2917.200 166.580 ;
        RECT 0.525 163.180 2917.600 164.580 ;
        RECT 2.800 161.180 2917.600 163.180 ;
        RECT 0.525 99.940 2917.600 161.180 ;
        RECT 0.525 97.940 2917.200 99.940 ;
        RECT 0.525 97.900 2917.600 97.940 ;
        RECT 2.800 95.900 2917.600 97.900 ;
        RECT 0.525 33.980 2917.600 95.900 ;
        RECT 0.525 33.300 2917.200 33.980 ;
        RECT 2.800 31.980 2917.200 33.300 ;
        RECT 2.800 31.300 2917.600 31.980 ;
        RECT 0.525 0.175 2917.600 31.300 ;
      LAYER met4 ;
        RECT 5.815 9.015 23.570 3512.705 ;
        RECT 27.470 9.015 55.820 3512.705 ;
        RECT 59.720 3442.745 88.070 3512.705 ;
        RECT 91.970 3442.745 120.320 3512.705 ;
        RECT 124.220 3442.745 152.570 3512.705 ;
        RECT 156.470 3442.745 184.820 3512.705 ;
        RECT 188.720 3442.745 217.070 3512.705 ;
        RECT 220.970 3442.745 249.320 3512.705 ;
        RECT 253.220 3442.745 281.570 3512.705 ;
        RECT 59.720 3226.400 281.570 3442.745 ;
        RECT 59.720 3166.745 88.070 3226.400 ;
        RECT 91.970 3166.745 120.320 3226.400 ;
        RECT 124.220 3166.745 152.570 3226.400 ;
        RECT 156.470 3166.745 184.820 3226.400 ;
        RECT 188.720 3166.745 217.070 3226.400 ;
        RECT 220.970 3166.745 249.320 3226.400 ;
        RECT 253.220 3166.745 281.570 3226.400 ;
        RECT 59.720 2950.400 281.570 3166.745 ;
        RECT 59.720 2890.745 88.070 2950.400 ;
        RECT 91.970 2890.745 120.320 2950.400 ;
        RECT 124.220 2890.745 152.570 2950.400 ;
        RECT 156.470 2890.745 184.820 2950.400 ;
        RECT 188.720 2890.745 217.070 2950.400 ;
        RECT 220.970 2890.745 249.320 2950.400 ;
        RECT 253.220 2890.745 281.570 2950.400 ;
        RECT 59.720 2674.400 281.570 2890.745 ;
        RECT 59.720 2614.745 88.070 2674.400 ;
        RECT 91.970 2614.745 120.320 2674.400 ;
        RECT 124.220 2614.745 152.570 2674.400 ;
        RECT 156.470 2614.745 184.820 2674.400 ;
        RECT 188.720 2614.745 217.070 2674.400 ;
        RECT 220.970 2614.745 249.320 2674.400 ;
        RECT 253.220 2614.745 281.570 2674.400 ;
        RECT 59.720 2398.400 281.570 2614.745 ;
        RECT 59.720 2338.745 88.070 2398.400 ;
        RECT 91.970 2338.745 120.320 2398.400 ;
        RECT 124.220 2338.745 152.570 2398.400 ;
        RECT 156.470 2338.745 184.820 2398.400 ;
        RECT 188.720 2338.745 217.070 2398.400 ;
        RECT 220.970 2338.745 249.320 2398.400 ;
        RECT 253.220 2338.745 281.570 2398.400 ;
        RECT 59.720 2122.400 281.570 2338.745 ;
        RECT 59.720 2062.745 88.070 2122.400 ;
        RECT 91.970 2062.745 120.320 2122.400 ;
        RECT 124.220 2062.745 152.570 2122.400 ;
        RECT 156.470 2062.745 184.820 2122.400 ;
        RECT 188.720 2062.745 217.070 2122.400 ;
        RECT 220.970 2062.745 249.320 2122.400 ;
        RECT 253.220 2062.745 281.570 2122.400 ;
        RECT 59.720 1846.400 281.570 2062.745 ;
        RECT 59.720 1786.745 88.070 1846.400 ;
        RECT 91.970 1786.745 120.320 1846.400 ;
        RECT 124.220 1786.745 152.570 1846.400 ;
        RECT 156.470 1786.745 184.820 1846.400 ;
        RECT 188.720 1786.745 217.070 1846.400 ;
        RECT 220.970 1786.745 249.320 1846.400 ;
        RECT 253.220 1786.745 281.570 1846.400 ;
        RECT 59.720 1570.400 281.570 1786.745 ;
        RECT 59.720 1510.745 88.070 1570.400 ;
        RECT 91.970 1510.745 120.320 1570.400 ;
        RECT 124.220 1510.745 152.570 1570.400 ;
        RECT 156.470 1510.745 184.820 1570.400 ;
        RECT 188.720 1510.745 217.070 1570.400 ;
        RECT 220.970 1510.745 249.320 1570.400 ;
        RECT 253.220 1510.745 281.570 1570.400 ;
        RECT 59.720 1294.400 281.570 1510.745 ;
        RECT 59.720 1234.745 88.070 1294.400 ;
        RECT 91.970 1234.745 120.320 1294.400 ;
        RECT 124.220 1234.745 152.570 1294.400 ;
        RECT 156.470 1234.745 184.820 1294.400 ;
        RECT 188.720 1234.745 217.070 1294.400 ;
        RECT 220.970 1234.745 249.320 1294.400 ;
        RECT 253.220 1234.745 281.570 1294.400 ;
        RECT 59.720 1018.400 281.570 1234.745 ;
        RECT 59.720 958.745 88.070 1018.400 ;
        RECT 91.970 958.745 120.320 1018.400 ;
        RECT 124.220 958.745 152.570 1018.400 ;
        RECT 156.470 958.745 184.820 1018.400 ;
        RECT 188.720 958.745 217.070 1018.400 ;
        RECT 220.970 958.745 249.320 1018.400 ;
        RECT 253.220 958.745 281.570 1018.400 ;
        RECT 59.720 742.400 281.570 958.745 ;
        RECT 59.720 682.745 88.070 742.400 ;
        RECT 91.970 682.745 120.320 742.400 ;
        RECT 124.220 682.745 152.570 742.400 ;
        RECT 156.470 682.745 184.820 742.400 ;
        RECT 188.720 682.745 217.070 742.400 ;
        RECT 220.970 682.745 249.320 742.400 ;
        RECT 253.220 682.745 281.570 742.400 ;
        RECT 59.720 466.400 281.570 682.745 ;
        RECT 59.720 406.745 88.070 466.400 ;
        RECT 91.970 406.745 120.320 466.400 ;
        RECT 124.220 406.745 152.570 466.400 ;
        RECT 156.470 406.745 184.820 466.400 ;
        RECT 188.720 406.745 217.070 466.400 ;
        RECT 220.970 406.745 249.320 466.400 ;
        RECT 253.220 406.745 281.570 466.400 ;
        RECT 59.720 190.400 281.570 406.745 ;
        RECT 59.720 9.015 88.070 190.400 ;
        RECT 91.970 9.015 120.320 190.400 ;
        RECT 124.220 9.015 152.570 190.400 ;
        RECT 156.470 9.015 184.820 190.400 ;
        RECT 188.720 9.015 217.070 190.400 ;
        RECT 220.970 9.015 249.320 190.400 ;
        RECT 253.220 9.015 281.570 190.400 ;
        RECT 285.470 9.015 313.820 3512.705 ;
        RECT 317.720 3442.745 346.070 3512.705 ;
        RECT 349.970 3442.745 378.320 3512.705 ;
        RECT 382.220 3442.745 410.570 3512.705 ;
        RECT 414.470 3442.745 442.820 3512.705 ;
        RECT 446.720 3442.745 475.070 3512.705 ;
        RECT 478.970 3442.745 507.320 3512.705 ;
        RECT 511.220 3442.745 539.570 3512.705 ;
        RECT 317.720 3226.400 539.570 3442.745 ;
        RECT 317.720 3166.745 346.070 3226.400 ;
        RECT 349.970 3166.745 378.320 3226.400 ;
        RECT 382.220 3166.745 410.570 3226.400 ;
        RECT 414.470 3166.745 442.820 3226.400 ;
        RECT 446.720 3166.745 475.070 3226.400 ;
        RECT 478.970 3166.745 507.320 3226.400 ;
        RECT 511.220 3166.745 539.570 3226.400 ;
        RECT 317.720 2950.400 539.570 3166.745 ;
        RECT 317.720 2890.745 346.070 2950.400 ;
        RECT 349.970 2890.745 378.320 2950.400 ;
        RECT 382.220 2890.745 410.570 2950.400 ;
        RECT 414.470 2890.745 442.820 2950.400 ;
        RECT 446.720 2890.745 475.070 2950.400 ;
        RECT 478.970 2890.745 507.320 2950.400 ;
        RECT 511.220 2890.745 539.570 2950.400 ;
        RECT 317.720 2674.400 539.570 2890.745 ;
        RECT 317.720 2614.745 346.070 2674.400 ;
        RECT 349.970 2614.745 378.320 2674.400 ;
        RECT 382.220 2614.745 410.570 2674.400 ;
        RECT 414.470 2614.745 442.820 2674.400 ;
        RECT 446.720 2614.745 475.070 2674.400 ;
        RECT 478.970 2614.745 507.320 2674.400 ;
        RECT 511.220 2614.745 539.570 2674.400 ;
        RECT 317.720 2398.400 539.570 2614.745 ;
        RECT 317.720 2338.745 346.070 2398.400 ;
        RECT 349.970 2338.745 378.320 2398.400 ;
        RECT 382.220 2338.745 410.570 2398.400 ;
        RECT 414.470 2338.745 442.820 2398.400 ;
        RECT 446.720 2338.745 475.070 2398.400 ;
        RECT 478.970 2338.745 507.320 2398.400 ;
        RECT 511.220 2338.745 539.570 2398.400 ;
        RECT 317.720 2122.400 539.570 2338.745 ;
        RECT 317.720 2062.745 346.070 2122.400 ;
        RECT 349.970 2062.745 378.320 2122.400 ;
        RECT 382.220 2062.745 410.570 2122.400 ;
        RECT 414.470 2062.745 442.820 2122.400 ;
        RECT 446.720 2062.745 475.070 2122.400 ;
        RECT 478.970 2062.745 507.320 2122.400 ;
        RECT 511.220 2062.745 539.570 2122.400 ;
        RECT 317.720 1846.400 539.570 2062.745 ;
        RECT 317.720 1786.745 346.070 1846.400 ;
        RECT 349.970 1786.745 378.320 1846.400 ;
        RECT 382.220 1786.745 410.570 1846.400 ;
        RECT 414.470 1786.745 442.820 1846.400 ;
        RECT 446.720 1786.745 475.070 1846.400 ;
        RECT 478.970 1786.745 507.320 1846.400 ;
        RECT 511.220 1786.745 539.570 1846.400 ;
        RECT 317.720 1570.400 539.570 1786.745 ;
        RECT 317.720 1510.745 346.070 1570.400 ;
        RECT 349.970 1510.745 378.320 1570.400 ;
        RECT 382.220 1510.745 410.570 1570.400 ;
        RECT 414.470 1510.745 442.820 1570.400 ;
        RECT 446.720 1510.745 475.070 1570.400 ;
        RECT 478.970 1510.745 507.320 1570.400 ;
        RECT 511.220 1510.745 539.570 1570.400 ;
        RECT 317.720 1294.400 539.570 1510.745 ;
        RECT 317.720 1234.745 346.070 1294.400 ;
        RECT 349.970 1234.745 378.320 1294.400 ;
        RECT 382.220 1234.745 410.570 1294.400 ;
        RECT 414.470 1234.745 442.820 1294.400 ;
        RECT 446.720 1234.745 475.070 1294.400 ;
        RECT 478.970 1234.745 507.320 1294.400 ;
        RECT 511.220 1234.745 539.570 1294.400 ;
        RECT 317.720 1018.400 539.570 1234.745 ;
        RECT 317.720 958.745 346.070 1018.400 ;
        RECT 349.970 958.745 378.320 1018.400 ;
        RECT 382.220 958.745 410.570 1018.400 ;
        RECT 414.470 958.745 442.820 1018.400 ;
        RECT 446.720 958.745 475.070 1018.400 ;
        RECT 478.970 958.745 507.320 1018.400 ;
        RECT 511.220 958.745 539.570 1018.400 ;
        RECT 317.720 742.400 539.570 958.745 ;
        RECT 317.720 682.745 346.070 742.400 ;
        RECT 349.970 682.745 378.320 742.400 ;
        RECT 382.220 682.745 410.570 742.400 ;
        RECT 414.470 682.745 442.820 742.400 ;
        RECT 446.720 682.745 475.070 742.400 ;
        RECT 478.970 682.745 507.320 742.400 ;
        RECT 511.220 682.745 539.570 742.400 ;
        RECT 317.720 466.400 539.570 682.745 ;
        RECT 317.720 406.745 346.070 466.400 ;
        RECT 349.970 406.745 378.320 466.400 ;
        RECT 382.220 406.745 410.570 466.400 ;
        RECT 414.470 406.745 442.820 466.400 ;
        RECT 446.720 406.745 475.070 466.400 ;
        RECT 478.970 406.745 507.320 466.400 ;
        RECT 511.220 406.745 539.570 466.400 ;
        RECT 317.720 190.400 539.570 406.745 ;
        RECT 317.720 9.015 346.070 190.400 ;
        RECT 349.970 9.015 378.320 190.400 ;
        RECT 382.220 9.015 410.570 190.400 ;
        RECT 414.470 9.015 442.820 190.400 ;
        RECT 446.720 9.015 475.070 190.400 ;
        RECT 478.970 9.015 507.320 190.400 ;
        RECT 511.220 9.015 539.570 190.400 ;
        RECT 543.470 9.015 571.820 3512.705 ;
        RECT 575.720 3442.745 604.070 3512.705 ;
        RECT 607.970 3442.745 636.320 3512.705 ;
        RECT 640.220 3442.745 668.570 3512.705 ;
        RECT 672.470 3442.745 700.820 3512.705 ;
        RECT 704.720 3442.745 733.070 3512.705 ;
        RECT 736.970 3442.745 765.320 3512.705 ;
        RECT 769.220 3442.745 797.570 3512.705 ;
        RECT 575.720 3226.400 797.570 3442.745 ;
        RECT 575.720 3166.745 604.070 3226.400 ;
        RECT 607.970 3166.745 636.320 3226.400 ;
        RECT 640.220 3166.745 668.570 3226.400 ;
        RECT 672.470 3166.745 700.820 3226.400 ;
        RECT 704.720 3166.745 733.070 3226.400 ;
        RECT 736.970 3166.745 765.320 3226.400 ;
        RECT 769.220 3166.745 797.570 3226.400 ;
        RECT 575.720 2950.400 797.570 3166.745 ;
        RECT 575.720 2890.745 604.070 2950.400 ;
        RECT 607.970 2890.745 636.320 2950.400 ;
        RECT 640.220 2890.745 668.570 2950.400 ;
        RECT 672.470 2890.745 700.820 2950.400 ;
        RECT 704.720 2890.745 733.070 2950.400 ;
        RECT 736.970 2890.745 765.320 2950.400 ;
        RECT 769.220 2890.745 797.570 2950.400 ;
        RECT 575.720 2674.400 797.570 2890.745 ;
        RECT 575.720 2614.745 604.070 2674.400 ;
        RECT 607.970 2614.745 636.320 2674.400 ;
        RECT 640.220 2614.745 668.570 2674.400 ;
        RECT 672.470 2614.745 700.820 2674.400 ;
        RECT 704.720 2614.745 733.070 2674.400 ;
        RECT 736.970 2614.745 765.320 2674.400 ;
        RECT 769.220 2614.745 797.570 2674.400 ;
        RECT 575.720 2398.400 797.570 2614.745 ;
        RECT 575.720 2338.745 604.070 2398.400 ;
        RECT 607.970 2338.745 636.320 2398.400 ;
        RECT 640.220 2338.745 668.570 2398.400 ;
        RECT 672.470 2338.745 700.820 2398.400 ;
        RECT 704.720 2338.745 733.070 2398.400 ;
        RECT 736.970 2338.745 765.320 2398.400 ;
        RECT 769.220 2338.745 797.570 2398.400 ;
        RECT 575.720 2122.400 797.570 2338.745 ;
        RECT 575.720 2062.745 604.070 2122.400 ;
        RECT 607.970 2062.745 636.320 2122.400 ;
        RECT 640.220 2062.745 668.570 2122.400 ;
        RECT 672.470 2062.745 700.820 2122.400 ;
        RECT 704.720 2062.745 733.070 2122.400 ;
        RECT 736.970 2062.745 765.320 2122.400 ;
        RECT 769.220 2062.745 797.570 2122.400 ;
        RECT 575.720 1846.400 797.570 2062.745 ;
        RECT 575.720 1786.745 604.070 1846.400 ;
        RECT 607.970 1786.745 636.320 1846.400 ;
        RECT 640.220 1786.745 668.570 1846.400 ;
        RECT 672.470 1786.745 700.820 1846.400 ;
        RECT 704.720 1786.745 733.070 1846.400 ;
        RECT 736.970 1786.745 765.320 1846.400 ;
        RECT 769.220 1786.745 797.570 1846.400 ;
        RECT 575.720 1570.400 797.570 1786.745 ;
        RECT 575.720 1510.745 604.070 1570.400 ;
        RECT 607.970 1510.745 636.320 1570.400 ;
        RECT 640.220 1510.745 668.570 1570.400 ;
        RECT 672.470 1510.745 700.820 1570.400 ;
        RECT 704.720 1510.745 733.070 1570.400 ;
        RECT 736.970 1510.745 765.320 1570.400 ;
        RECT 769.220 1510.745 797.570 1570.400 ;
        RECT 575.720 1294.400 797.570 1510.745 ;
        RECT 575.720 1234.745 604.070 1294.400 ;
        RECT 607.970 1234.745 636.320 1294.400 ;
        RECT 640.220 1234.745 668.570 1294.400 ;
        RECT 672.470 1234.745 700.820 1294.400 ;
        RECT 704.720 1234.745 733.070 1294.400 ;
        RECT 736.970 1234.745 765.320 1294.400 ;
        RECT 769.220 1234.745 797.570 1294.400 ;
        RECT 575.720 1018.400 797.570 1234.745 ;
        RECT 575.720 958.745 604.070 1018.400 ;
        RECT 607.970 958.745 636.320 1018.400 ;
        RECT 640.220 958.745 668.570 1018.400 ;
        RECT 672.470 958.745 700.820 1018.400 ;
        RECT 704.720 958.745 733.070 1018.400 ;
        RECT 736.970 958.745 765.320 1018.400 ;
        RECT 769.220 958.745 797.570 1018.400 ;
        RECT 575.720 742.400 797.570 958.745 ;
        RECT 575.720 682.745 604.070 742.400 ;
        RECT 607.970 682.745 636.320 742.400 ;
        RECT 640.220 682.745 668.570 742.400 ;
        RECT 672.470 682.745 700.820 742.400 ;
        RECT 704.720 682.745 733.070 742.400 ;
        RECT 736.970 682.745 765.320 742.400 ;
        RECT 769.220 682.745 797.570 742.400 ;
        RECT 575.720 466.400 797.570 682.745 ;
        RECT 575.720 406.745 604.070 466.400 ;
        RECT 607.970 406.745 636.320 466.400 ;
        RECT 640.220 406.745 668.570 466.400 ;
        RECT 672.470 406.745 700.820 466.400 ;
        RECT 704.720 406.745 733.070 466.400 ;
        RECT 736.970 406.745 765.320 466.400 ;
        RECT 769.220 406.745 797.570 466.400 ;
        RECT 575.720 190.400 797.570 406.745 ;
        RECT 575.720 9.015 604.070 190.400 ;
        RECT 607.970 9.015 636.320 190.400 ;
        RECT 640.220 9.015 668.570 190.400 ;
        RECT 672.470 9.015 700.820 190.400 ;
        RECT 704.720 9.015 733.070 190.400 ;
        RECT 736.970 9.015 765.320 190.400 ;
        RECT 769.220 9.015 797.570 190.400 ;
        RECT 801.470 9.015 829.820 3512.705 ;
        RECT 833.720 3442.745 862.070 3512.705 ;
        RECT 865.970 3442.745 894.320 3512.705 ;
        RECT 898.220 3442.745 926.570 3512.705 ;
        RECT 930.470 3442.745 958.820 3512.705 ;
        RECT 962.720 3442.745 991.070 3512.705 ;
        RECT 994.970 3442.745 1023.320 3512.705 ;
        RECT 1027.220 3442.745 1055.570 3512.705 ;
        RECT 833.720 3226.400 1055.570 3442.745 ;
        RECT 833.720 3166.745 862.070 3226.400 ;
        RECT 865.970 3166.745 894.320 3226.400 ;
        RECT 898.220 3166.745 926.570 3226.400 ;
        RECT 930.470 3166.745 958.820 3226.400 ;
        RECT 962.720 3166.745 991.070 3226.400 ;
        RECT 994.970 3166.745 1023.320 3226.400 ;
        RECT 1027.220 3166.745 1055.570 3226.400 ;
        RECT 833.720 2950.400 1055.570 3166.745 ;
        RECT 833.720 2890.745 862.070 2950.400 ;
        RECT 865.970 2890.745 894.320 2950.400 ;
        RECT 898.220 2890.745 926.570 2950.400 ;
        RECT 930.470 2890.745 958.820 2950.400 ;
        RECT 962.720 2890.745 991.070 2950.400 ;
        RECT 994.970 2890.745 1023.320 2950.400 ;
        RECT 1027.220 2890.745 1055.570 2950.400 ;
        RECT 833.720 2674.400 1055.570 2890.745 ;
        RECT 833.720 2614.745 862.070 2674.400 ;
        RECT 865.970 2614.745 894.320 2674.400 ;
        RECT 898.220 2614.745 926.570 2674.400 ;
        RECT 930.470 2614.745 958.820 2674.400 ;
        RECT 962.720 2614.745 991.070 2674.400 ;
        RECT 994.970 2614.745 1023.320 2674.400 ;
        RECT 1027.220 2614.745 1055.570 2674.400 ;
        RECT 833.720 2398.400 1055.570 2614.745 ;
        RECT 833.720 2338.745 862.070 2398.400 ;
        RECT 865.970 2338.745 894.320 2398.400 ;
        RECT 898.220 2338.745 926.570 2398.400 ;
        RECT 930.470 2338.745 958.820 2398.400 ;
        RECT 962.720 2338.745 991.070 2398.400 ;
        RECT 994.970 2338.745 1023.320 2398.400 ;
        RECT 1027.220 2338.745 1055.570 2398.400 ;
        RECT 833.720 2122.400 1055.570 2338.745 ;
        RECT 833.720 2062.745 862.070 2122.400 ;
        RECT 865.970 2062.745 894.320 2122.400 ;
        RECT 898.220 2062.745 926.570 2122.400 ;
        RECT 930.470 2062.745 958.820 2122.400 ;
        RECT 962.720 2062.745 991.070 2122.400 ;
        RECT 994.970 2062.745 1023.320 2122.400 ;
        RECT 1027.220 2062.745 1055.570 2122.400 ;
        RECT 833.720 1846.400 1055.570 2062.745 ;
        RECT 833.720 1786.745 862.070 1846.400 ;
        RECT 865.970 1786.745 894.320 1846.400 ;
        RECT 898.220 1786.745 926.570 1846.400 ;
        RECT 930.470 1786.745 958.820 1846.400 ;
        RECT 962.720 1786.745 991.070 1846.400 ;
        RECT 994.970 1786.745 1023.320 1846.400 ;
        RECT 1027.220 1786.745 1055.570 1846.400 ;
        RECT 833.720 1570.400 1055.570 1786.745 ;
        RECT 833.720 1510.745 862.070 1570.400 ;
        RECT 865.970 1510.745 894.320 1570.400 ;
        RECT 898.220 1510.745 926.570 1570.400 ;
        RECT 930.470 1510.745 958.820 1570.400 ;
        RECT 962.720 1510.745 991.070 1570.400 ;
        RECT 994.970 1510.745 1023.320 1570.400 ;
        RECT 1027.220 1510.745 1055.570 1570.400 ;
        RECT 833.720 1294.400 1055.570 1510.745 ;
        RECT 833.720 1234.745 862.070 1294.400 ;
        RECT 865.970 1234.745 894.320 1294.400 ;
        RECT 898.220 1234.745 926.570 1294.400 ;
        RECT 930.470 1234.745 958.820 1294.400 ;
        RECT 962.720 1234.745 991.070 1294.400 ;
        RECT 994.970 1234.745 1023.320 1294.400 ;
        RECT 1027.220 1234.745 1055.570 1294.400 ;
        RECT 833.720 1018.400 1055.570 1234.745 ;
        RECT 833.720 958.745 862.070 1018.400 ;
        RECT 865.970 958.745 894.320 1018.400 ;
        RECT 898.220 958.745 926.570 1018.400 ;
        RECT 930.470 958.745 958.820 1018.400 ;
        RECT 962.720 958.745 991.070 1018.400 ;
        RECT 994.970 958.745 1023.320 1018.400 ;
        RECT 1027.220 958.745 1055.570 1018.400 ;
        RECT 833.720 742.400 1055.570 958.745 ;
        RECT 833.720 682.745 862.070 742.400 ;
        RECT 865.970 682.745 894.320 742.400 ;
        RECT 898.220 682.745 926.570 742.400 ;
        RECT 930.470 682.745 958.820 742.400 ;
        RECT 962.720 682.745 991.070 742.400 ;
        RECT 994.970 682.745 1023.320 742.400 ;
        RECT 1027.220 682.745 1055.570 742.400 ;
        RECT 833.720 466.400 1055.570 682.745 ;
        RECT 833.720 406.745 862.070 466.400 ;
        RECT 865.970 406.745 894.320 466.400 ;
        RECT 898.220 406.745 926.570 466.400 ;
        RECT 930.470 406.745 958.820 466.400 ;
        RECT 962.720 406.745 991.070 466.400 ;
        RECT 994.970 406.745 1023.320 466.400 ;
        RECT 1027.220 406.745 1055.570 466.400 ;
        RECT 833.720 190.400 1055.570 406.745 ;
        RECT 833.720 9.015 862.070 190.400 ;
        RECT 865.970 9.015 894.320 190.400 ;
        RECT 898.220 9.015 926.570 190.400 ;
        RECT 930.470 9.015 958.820 190.400 ;
        RECT 962.720 9.015 991.070 190.400 ;
        RECT 994.970 9.015 1023.320 190.400 ;
        RECT 1027.220 9.015 1055.570 190.400 ;
        RECT 1059.470 9.015 1087.820 3512.705 ;
        RECT 1091.720 3442.745 1120.070 3512.705 ;
        RECT 1123.970 3442.745 1152.320 3512.705 ;
        RECT 1156.220 3442.745 1184.570 3512.705 ;
        RECT 1188.470 3442.745 1216.820 3512.705 ;
        RECT 1220.720 3442.745 1249.070 3512.705 ;
        RECT 1252.970 3442.745 1281.320 3512.705 ;
        RECT 1285.220 3442.745 1313.570 3512.705 ;
        RECT 1091.720 3226.400 1313.570 3442.745 ;
        RECT 1091.720 3166.745 1120.070 3226.400 ;
        RECT 1123.970 3166.745 1152.320 3226.400 ;
        RECT 1156.220 3166.745 1184.570 3226.400 ;
        RECT 1188.470 3166.745 1216.820 3226.400 ;
        RECT 1220.720 3166.745 1249.070 3226.400 ;
        RECT 1252.970 3166.745 1281.320 3226.400 ;
        RECT 1285.220 3166.745 1313.570 3226.400 ;
        RECT 1091.720 2950.400 1313.570 3166.745 ;
        RECT 1091.720 2890.745 1120.070 2950.400 ;
        RECT 1123.970 2890.745 1152.320 2950.400 ;
        RECT 1156.220 2890.745 1184.570 2950.400 ;
        RECT 1188.470 2890.745 1216.820 2950.400 ;
        RECT 1220.720 2890.745 1249.070 2950.400 ;
        RECT 1252.970 2890.745 1281.320 2950.400 ;
        RECT 1285.220 2890.745 1313.570 2950.400 ;
        RECT 1091.720 2674.400 1313.570 2890.745 ;
        RECT 1091.720 2614.745 1120.070 2674.400 ;
        RECT 1123.970 2614.745 1152.320 2674.400 ;
        RECT 1156.220 2614.745 1184.570 2674.400 ;
        RECT 1188.470 2614.745 1216.820 2674.400 ;
        RECT 1220.720 2614.745 1249.070 2674.400 ;
        RECT 1252.970 2614.745 1281.320 2674.400 ;
        RECT 1285.220 2614.745 1313.570 2674.400 ;
        RECT 1091.720 2398.400 1313.570 2614.745 ;
        RECT 1091.720 2338.745 1120.070 2398.400 ;
        RECT 1123.970 2338.745 1152.320 2398.400 ;
        RECT 1156.220 2338.745 1184.570 2398.400 ;
        RECT 1188.470 2338.745 1216.820 2398.400 ;
        RECT 1220.720 2338.745 1249.070 2398.400 ;
        RECT 1252.970 2338.745 1281.320 2398.400 ;
        RECT 1285.220 2338.745 1313.570 2398.400 ;
        RECT 1091.720 2122.400 1313.570 2338.745 ;
        RECT 1091.720 2062.745 1120.070 2122.400 ;
        RECT 1123.970 2062.745 1152.320 2122.400 ;
        RECT 1156.220 2062.745 1184.570 2122.400 ;
        RECT 1188.470 2062.745 1216.820 2122.400 ;
        RECT 1220.720 2062.745 1249.070 2122.400 ;
        RECT 1252.970 2062.745 1281.320 2122.400 ;
        RECT 1285.220 2062.745 1313.570 2122.400 ;
        RECT 1091.720 1846.400 1313.570 2062.745 ;
        RECT 1091.720 1786.745 1120.070 1846.400 ;
        RECT 1123.970 1786.745 1152.320 1846.400 ;
        RECT 1156.220 1786.745 1184.570 1846.400 ;
        RECT 1188.470 1786.745 1216.820 1846.400 ;
        RECT 1220.720 1786.745 1249.070 1846.400 ;
        RECT 1252.970 1786.745 1281.320 1846.400 ;
        RECT 1285.220 1786.745 1313.570 1846.400 ;
        RECT 1091.720 1570.400 1313.570 1786.745 ;
        RECT 1091.720 1510.745 1120.070 1570.400 ;
        RECT 1123.970 1510.745 1152.320 1570.400 ;
        RECT 1156.220 1510.745 1184.570 1570.400 ;
        RECT 1188.470 1510.745 1216.820 1570.400 ;
        RECT 1220.720 1510.745 1249.070 1570.400 ;
        RECT 1252.970 1510.745 1281.320 1570.400 ;
        RECT 1285.220 1510.745 1313.570 1570.400 ;
        RECT 1091.720 1294.400 1313.570 1510.745 ;
        RECT 1091.720 1234.745 1120.070 1294.400 ;
        RECT 1123.970 1234.745 1152.320 1294.400 ;
        RECT 1156.220 1234.745 1184.570 1294.400 ;
        RECT 1188.470 1234.745 1216.820 1294.400 ;
        RECT 1220.720 1234.745 1249.070 1294.400 ;
        RECT 1252.970 1234.745 1281.320 1294.400 ;
        RECT 1285.220 1234.745 1313.570 1294.400 ;
        RECT 1091.720 1018.400 1313.570 1234.745 ;
        RECT 1091.720 958.745 1120.070 1018.400 ;
        RECT 1123.970 958.745 1152.320 1018.400 ;
        RECT 1156.220 958.745 1184.570 1018.400 ;
        RECT 1188.470 958.745 1216.820 1018.400 ;
        RECT 1220.720 958.745 1249.070 1018.400 ;
        RECT 1252.970 958.745 1281.320 1018.400 ;
        RECT 1285.220 958.745 1313.570 1018.400 ;
        RECT 1091.720 742.400 1313.570 958.745 ;
        RECT 1091.720 682.745 1120.070 742.400 ;
        RECT 1123.970 682.745 1152.320 742.400 ;
        RECT 1156.220 682.745 1184.570 742.400 ;
        RECT 1188.470 682.745 1216.820 742.400 ;
        RECT 1220.720 682.745 1249.070 742.400 ;
        RECT 1252.970 682.745 1281.320 742.400 ;
        RECT 1285.220 682.745 1313.570 742.400 ;
        RECT 1091.720 466.400 1313.570 682.745 ;
        RECT 1091.720 406.745 1120.070 466.400 ;
        RECT 1123.970 406.745 1152.320 466.400 ;
        RECT 1156.220 406.745 1184.570 466.400 ;
        RECT 1188.470 406.745 1216.820 466.400 ;
        RECT 1220.720 406.745 1249.070 466.400 ;
        RECT 1252.970 406.745 1281.320 466.400 ;
        RECT 1285.220 406.745 1313.570 466.400 ;
        RECT 1091.720 190.400 1313.570 406.745 ;
        RECT 1091.720 9.015 1120.070 190.400 ;
        RECT 1123.970 9.015 1152.320 190.400 ;
        RECT 1156.220 9.015 1184.570 190.400 ;
        RECT 1188.470 9.015 1216.820 190.400 ;
        RECT 1220.720 9.015 1249.070 190.400 ;
        RECT 1252.970 9.015 1281.320 190.400 ;
        RECT 1285.220 9.015 1313.570 190.400 ;
        RECT 1317.470 9.015 1345.820 3512.705 ;
        RECT 1349.720 3442.745 1378.070 3512.705 ;
        RECT 1381.970 3442.745 1410.320 3512.705 ;
        RECT 1414.220 3442.745 1442.570 3512.705 ;
        RECT 1446.470 3442.745 1474.820 3512.705 ;
        RECT 1478.720 3442.745 1507.070 3512.705 ;
        RECT 1510.970 3442.745 1539.320 3512.705 ;
        RECT 1543.220 3442.745 1571.570 3512.705 ;
        RECT 1349.720 3226.400 1571.570 3442.745 ;
        RECT 1349.720 3166.745 1378.070 3226.400 ;
        RECT 1381.970 3166.745 1410.320 3226.400 ;
        RECT 1414.220 3166.745 1442.570 3226.400 ;
        RECT 1446.470 3166.745 1474.820 3226.400 ;
        RECT 1478.720 3166.745 1507.070 3226.400 ;
        RECT 1510.970 3166.745 1539.320 3226.400 ;
        RECT 1543.220 3166.745 1571.570 3226.400 ;
        RECT 1349.720 2950.400 1571.570 3166.745 ;
        RECT 1349.720 2890.745 1378.070 2950.400 ;
        RECT 1381.970 2890.745 1410.320 2950.400 ;
        RECT 1414.220 2890.745 1442.570 2950.400 ;
        RECT 1446.470 2890.745 1474.820 2950.400 ;
        RECT 1478.720 2890.745 1507.070 2950.400 ;
        RECT 1510.970 2890.745 1539.320 2950.400 ;
        RECT 1543.220 2890.745 1571.570 2950.400 ;
        RECT 1349.720 2674.400 1571.570 2890.745 ;
        RECT 1349.720 2614.745 1378.070 2674.400 ;
        RECT 1381.970 2614.745 1410.320 2674.400 ;
        RECT 1414.220 2614.745 1442.570 2674.400 ;
        RECT 1446.470 2614.745 1474.820 2674.400 ;
        RECT 1478.720 2614.745 1507.070 2674.400 ;
        RECT 1510.970 2614.745 1539.320 2674.400 ;
        RECT 1543.220 2614.745 1571.570 2674.400 ;
        RECT 1349.720 2398.400 1571.570 2614.745 ;
        RECT 1349.720 2338.745 1378.070 2398.400 ;
        RECT 1381.970 2338.745 1410.320 2398.400 ;
        RECT 1414.220 2338.745 1442.570 2398.400 ;
        RECT 1446.470 2338.745 1474.820 2398.400 ;
        RECT 1478.720 2338.745 1507.070 2398.400 ;
        RECT 1510.970 2338.745 1539.320 2398.400 ;
        RECT 1543.220 2338.745 1571.570 2398.400 ;
        RECT 1349.720 2122.400 1571.570 2338.745 ;
        RECT 1349.720 2062.745 1378.070 2122.400 ;
        RECT 1381.970 2062.745 1410.320 2122.400 ;
        RECT 1414.220 2062.745 1442.570 2122.400 ;
        RECT 1446.470 2062.745 1474.820 2122.400 ;
        RECT 1478.720 2062.745 1507.070 2122.400 ;
        RECT 1510.970 2062.745 1539.320 2122.400 ;
        RECT 1543.220 2062.745 1571.570 2122.400 ;
        RECT 1349.720 1846.400 1571.570 2062.745 ;
        RECT 1349.720 1786.745 1378.070 1846.400 ;
        RECT 1381.970 1786.745 1410.320 1846.400 ;
        RECT 1414.220 1786.745 1442.570 1846.400 ;
        RECT 1446.470 1786.745 1474.820 1846.400 ;
        RECT 1478.720 1786.745 1507.070 1846.400 ;
        RECT 1510.970 1786.745 1539.320 1846.400 ;
        RECT 1543.220 1786.745 1571.570 1846.400 ;
        RECT 1349.720 1570.400 1571.570 1786.745 ;
        RECT 1349.720 1510.745 1378.070 1570.400 ;
        RECT 1381.970 1510.745 1410.320 1570.400 ;
        RECT 1414.220 1510.745 1442.570 1570.400 ;
        RECT 1446.470 1510.745 1474.820 1570.400 ;
        RECT 1478.720 1510.745 1507.070 1570.400 ;
        RECT 1510.970 1510.745 1539.320 1570.400 ;
        RECT 1543.220 1510.745 1571.570 1570.400 ;
        RECT 1349.720 1294.400 1571.570 1510.745 ;
        RECT 1349.720 1234.745 1378.070 1294.400 ;
        RECT 1381.970 1234.745 1410.320 1294.400 ;
        RECT 1414.220 1234.745 1442.570 1294.400 ;
        RECT 1446.470 1234.745 1474.820 1294.400 ;
        RECT 1478.720 1234.745 1507.070 1294.400 ;
        RECT 1510.970 1234.745 1539.320 1294.400 ;
        RECT 1543.220 1234.745 1571.570 1294.400 ;
        RECT 1349.720 1018.400 1571.570 1234.745 ;
        RECT 1349.720 958.745 1378.070 1018.400 ;
        RECT 1381.970 958.745 1410.320 1018.400 ;
        RECT 1414.220 958.745 1442.570 1018.400 ;
        RECT 1446.470 958.745 1474.820 1018.400 ;
        RECT 1478.720 958.745 1507.070 1018.400 ;
        RECT 1510.970 958.745 1539.320 1018.400 ;
        RECT 1543.220 958.745 1571.570 1018.400 ;
        RECT 1349.720 742.400 1571.570 958.745 ;
        RECT 1349.720 682.745 1378.070 742.400 ;
        RECT 1381.970 682.745 1410.320 742.400 ;
        RECT 1414.220 682.745 1442.570 742.400 ;
        RECT 1446.470 682.745 1474.820 742.400 ;
        RECT 1478.720 682.745 1507.070 742.400 ;
        RECT 1510.970 682.745 1539.320 742.400 ;
        RECT 1543.220 682.745 1571.570 742.400 ;
        RECT 1349.720 466.400 1571.570 682.745 ;
        RECT 1349.720 406.745 1378.070 466.400 ;
        RECT 1381.970 406.745 1410.320 466.400 ;
        RECT 1414.220 406.745 1442.570 466.400 ;
        RECT 1446.470 406.745 1474.820 466.400 ;
        RECT 1478.720 406.745 1507.070 466.400 ;
        RECT 1510.970 406.745 1539.320 466.400 ;
        RECT 1543.220 406.745 1571.570 466.400 ;
        RECT 1349.720 190.400 1571.570 406.745 ;
        RECT 1349.720 9.015 1378.070 190.400 ;
        RECT 1381.970 9.015 1410.320 190.400 ;
        RECT 1414.220 9.015 1442.570 190.400 ;
        RECT 1446.470 9.015 1474.820 190.400 ;
        RECT 1478.720 9.015 1507.070 190.400 ;
        RECT 1510.970 9.015 1539.320 190.400 ;
        RECT 1543.220 9.015 1571.570 190.400 ;
        RECT 1575.470 9.015 1603.820 3512.705 ;
        RECT 1607.720 3442.745 1636.070 3512.705 ;
        RECT 1639.970 3442.745 1668.320 3512.705 ;
        RECT 1672.220 3442.745 1700.570 3512.705 ;
        RECT 1704.470 3442.745 1732.820 3512.705 ;
        RECT 1736.720 3442.745 1765.070 3512.705 ;
        RECT 1768.970 3442.745 1797.320 3512.705 ;
        RECT 1801.220 3442.745 1829.570 3512.705 ;
        RECT 1607.720 3226.400 1829.570 3442.745 ;
        RECT 1607.720 3166.745 1636.070 3226.400 ;
        RECT 1639.970 3166.745 1668.320 3226.400 ;
        RECT 1672.220 3166.745 1700.570 3226.400 ;
        RECT 1704.470 3166.745 1732.820 3226.400 ;
        RECT 1736.720 3166.745 1765.070 3226.400 ;
        RECT 1768.970 3166.745 1797.320 3226.400 ;
        RECT 1801.220 3166.745 1829.570 3226.400 ;
        RECT 1607.720 2950.400 1829.570 3166.745 ;
        RECT 1607.720 2890.745 1636.070 2950.400 ;
        RECT 1639.970 2890.745 1668.320 2950.400 ;
        RECT 1672.220 2890.745 1700.570 2950.400 ;
        RECT 1704.470 2890.745 1732.820 2950.400 ;
        RECT 1736.720 2890.745 1765.070 2950.400 ;
        RECT 1768.970 2890.745 1797.320 2950.400 ;
        RECT 1801.220 2890.745 1829.570 2950.400 ;
        RECT 1607.720 2674.400 1829.570 2890.745 ;
        RECT 1607.720 2614.745 1636.070 2674.400 ;
        RECT 1639.970 2614.745 1668.320 2674.400 ;
        RECT 1672.220 2614.745 1700.570 2674.400 ;
        RECT 1704.470 2614.745 1732.820 2674.400 ;
        RECT 1736.720 2614.745 1765.070 2674.400 ;
        RECT 1768.970 2614.745 1797.320 2674.400 ;
        RECT 1801.220 2614.745 1829.570 2674.400 ;
        RECT 1607.720 2398.400 1829.570 2614.745 ;
        RECT 1607.720 2338.745 1636.070 2398.400 ;
        RECT 1639.970 2338.745 1668.320 2398.400 ;
        RECT 1672.220 2338.745 1700.570 2398.400 ;
        RECT 1704.470 2338.745 1732.820 2398.400 ;
        RECT 1736.720 2338.745 1765.070 2398.400 ;
        RECT 1768.970 2338.745 1797.320 2398.400 ;
        RECT 1801.220 2338.745 1829.570 2398.400 ;
        RECT 1607.720 2122.400 1829.570 2338.745 ;
        RECT 1607.720 2062.745 1636.070 2122.400 ;
        RECT 1639.970 2062.745 1668.320 2122.400 ;
        RECT 1672.220 2062.745 1700.570 2122.400 ;
        RECT 1704.470 2062.745 1732.820 2122.400 ;
        RECT 1736.720 2062.745 1765.070 2122.400 ;
        RECT 1768.970 2062.745 1797.320 2122.400 ;
        RECT 1801.220 2062.745 1829.570 2122.400 ;
        RECT 1607.720 1846.400 1829.570 2062.745 ;
        RECT 1607.720 1786.745 1636.070 1846.400 ;
        RECT 1639.970 1786.745 1668.320 1846.400 ;
        RECT 1672.220 1786.745 1700.570 1846.400 ;
        RECT 1704.470 1786.745 1732.820 1846.400 ;
        RECT 1736.720 1786.745 1765.070 1846.400 ;
        RECT 1768.970 1786.745 1797.320 1846.400 ;
        RECT 1801.220 1786.745 1829.570 1846.400 ;
        RECT 1607.720 1570.400 1829.570 1786.745 ;
        RECT 1607.720 1510.745 1636.070 1570.400 ;
        RECT 1639.970 1510.745 1668.320 1570.400 ;
        RECT 1672.220 1510.745 1700.570 1570.400 ;
        RECT 1704.470 1510.745 1732.820 1570.400 ;
        RECT 1736.720 1510.745 1765.070 1570.400 ;
        RECT 1768.970 1510.745 1797.320 1570.400 ;
        RECT 1801.220 1510.745 1829.570 1570.400 ;
        RECT 1607.720 1294.400 1829.570 1510.745 ;
        RECT 1607.720 1234.745 1636.070 1294.400 ;
        RECT 1639.970 1234.745 1668.320 1294.400 ;
        RECT 1672.220 1234.745 1700.570 1294.400 ;
        RECT 1704.470 1234.745 1732.820 1294.400 ;
        RECT 1736.720 1234.745 1765.070 1294.400 ;
        RECT 1768.970 1234.745 1797.320 1294.400 ;
        RECT 1801.220 1234.745 1829.570 1294.400 ;
        RECT 1607.720 1018.400 1829.570 1234.745 ;
        RECT 1607.720 958.745 1636.070 1018.400 ;
        RECT 1639.970 958.745 1668.320 1018.400 ;
        RECT 1672.220 958.745 1700.570 1018.400 ;
        RECT 1704.470 958.745 1732.820 1018.400 ;
        RECT 1736.720 958.745 1765.070 1018.400 ;
        RECT 1768.970 958.745 1797.320 1018.400 ;
        RECT 1801.220 958.745 1829.570 1018.400 ;
        RECT 1607.720 742.400 1829.570 958.745 ;
        RECT 1607.720 682.745 1636.070 742.400 ;
        RECT 1639.970 682.745 1668.320 742.400 ;
        RECT 1672.220 682.745 1700.570 742.400 ;
        RECT 1704.470 682.745 1732.820 742.400 ;
        RECT 1736.720 682.745 1765.070 742.400 ;
        RECT 1768.970 682.745 1797.320 742.400 ;
        RECT 1801.220 682.745 1829.570 742.400 ;
        RECT 1607.720 466.400 1829.570 682.745 ;
        RECT 1607.720 406.745 1636.070 466.400 ;
        RECT 1639.970 406.745 1668.320 466.400 ;
        RECT 1672.220 406.745 1700.570 466.400 ;
        RECT 1704.470 406.745 1732.820 466.400 ;
        RECT 1736.720 406.745 1765.070 466.400 ;
        RECT 1768.970 406.745 1797.320 466.400 ;
        RECT 1801.220 406.745 1829.570 466.400 ;
        RECT 1607.720 190.400 1829.570 406.745 ;
        RECT 1607.720 9.015 1636.070 190.400 ;
        RECT 1639.970 9.015 1668.320 190.400 ;
        RECT 1672.220 9.015 1700.570 190.400 ;
        RECT 1704.470 9.015 1732.820 190.400 ;
        RECT 1736.720 9.015 1765.070 190.400 ;
        RECT 1768.970 9.015 1797.320 190.400 ;
        RECT 1801.220 9.015 1829.570 190.400 ;
        RECT 1833.470 9.015 1861.820 3512.705 ;
        RECT 1865.720 3442.745 1894.070 3512.705 ;
        RECT 1897.970 3442.745 1926.320 3512.705 ;
        RECT 1930.220 3442.745 1958.570 3512.705 ;
        RECT 1962.470 3442.745 1990.820 3512.705 ;
        RECT 1994.720 3442.745 2023.070 3512.705 ;
        RECT 2026.970 3442.745 2055.320 3512.705 ;
        RECT 2059.220 3442.745 2087.570 3512.705 ;
        RECT 1865.720 3226.400 2087.570 3442.745 ;
        RECT 1865.720 3166.745 1894.070 3226.400 ;
        RECT 1897.970 3166.745 1926.320 3226.400 ;
        RECT 1930.220 3166.745 1958.570 3226.400 ;
        RECT 1962.470 3166.745 1990.820 3226.400 ;
        RECT 1994.720 3166.745 2023.070 3226.400 ;
        RECT 2026.970 3166.745 2055.320 3226.400 ;
        RECT 2059.220 3166.745 2087.570 3226.400 ;
        RECT 1865.720 2950.400 2087.570 3166.745 ;
        RECT 1865.720 2890.745 1894.070 2950.400 ;
        RECT 1897.970 2890.745 1926.320 2950.400 ;
        RECT 1930.220 2890.745 1958.570 2950.400 ;
        RECT 1962.470 2890.745 1990.820 2950.400 ;
        RECT 1994.720 2890.745 2023.070 2950.400 ;
        RECT 2026.970 2890.745 2055.320 2950.400 ;
        RECT 2059.220 2890.745 2087.570 2950.400 ;
        RECT 1865.720 2674.400 2087.570 2890.745 ;
        RECT 1865.720 2614.745 1894.070 2674.400 ;
        RECT 1897.970 2614.745 1926.320 2674.400 ;
        RECT 1930.220 2614.745 1958.570 2674.400 ;
        RECT 1962.470 2614.745 1990.820 2674.400 ;
        RECT 1994.720 2614.745 2023.070 2674.400 ;
        RECT 2026.970 2614.745 2055.320 2674.400 ;
        RECT 2059.220 2614.745 2087.570 2674.400 ;
        RECT 1865.720 2398.400 2087.570 2614.745 ;
        RECT 1865.720 2338.745 1894.070 2398.400 ;
        RECT 1897.970 2338.745 1926.320 2398.400 ;
        RECT 1930.220 2338.745 1958.570 2398.400 ;
        RECT 1962.470 2338.745 1990.820 2398.400 ;
        RECT 1994.720 2338.745 2023.070 2398.400 ;
        RECT 2026.970 2338.745 2055.320 2398.400 ;
        RECT 2059.220 2338.745 2087.570 2398.400 ;
        RECT 1865.720 2122.400 2087.570 2338.745 ;
        RECT 1865.720 2062.745 1894.070 2122.400 ;
        RECT 1897.970 2062.745 1926.320 2122.400 ;
        RECT 1930.220 2062.745 1958.570 2122.400 ;
        RECT 1962.470 2062.745 1990.820 2122.400 ;
        RECT 1994.720 2062.745 2023.070 2122.400 ;
        RECT 2026.970 2062.745 2055.320 2122.400 ;
        RECT 2059.220 2062.745 2087.570 2122.400 ;
        RECT 1865.720 1846.400 2087.570 2062.745 ;
        RECT 1865.720 1786.745 1894.070 1846.400 ;
        RECT 1897.970 1786.745 1926.320 1846.400 ;
        RECT 1930.220 1786.745 1958.570 1846.400 ;
        RECT 1962.470 1786.745 1990.820 1846.400 ;
        RECT 1994.720 1786.745 2023.070 1846.400 ;
        RECT 2026.970 1786.745 2055.320 1846.400 ;
        RECT 2059.220 1786.745 2087.570 1846.400 ;
        RECT 1865.720 1570.400 2087.570 1786.745 ;
        RECT 1865.720 1510.745 1894.070 1570.400 ;
        RECT 1897.970 1510.745 1926.320 1570.400 ;
        RECT 1930.220 1510.745 1958.570 1570.400 ;
        RECT 1962.470 1510.745 1990.820 1570.400 ;
        RECT 1994.720 1510.745 2023.070 1570.400 ;
        RECT 2026.970 1510.745 2055.320 1570.400 ;
        RECT 2059.220 1510.745 2087.570 1570.400 ;
        RECT 1865.720 1294.400 2087.570 1510.745 ;
        RECT 1865.720 1234.745 1894.070 1294.400 ;
        RECT 1897.970 1234.745 1926.320 1294.400 ;
        RECT 1930.220 1234.745 1958.570 1294.400 ;
        RECT 1962.470 1234.745 1990.820 1294.400 ;
        RECT 1994.720 1234.745 2023.070 1294.400 ;
        RECT 2026.970 1234.745 2055.320 1294.400 ;
        RECT 2059.220 1234.745 2087.570 1294.400 ;
        RECT 1865.720 1018.400 2087.570 1234.745 ;
        RECT 1865.720 958.745 1894.070 1018.400 ;
        RECT 1897.970 958.745 1926.320 1018.400 ;
        RECT 1930.220 958.745 1958.570 1018.400 ;
        RECT 1962.470 958.745 1990.820 1018.400 ;
        RECT 1994.720 958.745 2023.070 1018.400 ;
        RECT 2026.970 958.745 2055.320 1018.400 ;
        RECT 2059.220 958.745 2087.570 1018.400 ;
        RECT 1865.720 742.400 2087.570 958.745 ;
        RECT 1865.720 682.745 1894.070 742.400 ;
        RECT 1897.970 682.745 1926.320 742.400 ;
        RECT 1930.220 682.745 1958.570 742.400 ;
        RECT 1962.470 682.745 1990.820 742.400 ;
        RECT 1994.720 682.745 2023.070 742.400 ;
        RECT 2026.970 682.745 2055.320 742.400 ;
        RECT 2059.220 682.745 2087.570 742.400 ;
        RECT 1865.720 466.400 2087.570 682.745 ;
        RECT 1865.720 406.745 1894.070 466.400 ;
        RECT 1897.970 406.745 1926.320 466.400 ;
        RECT 1930.220 406.745 1958.570 466.400 ;
        RECT 1962.470 406.745 1990.820 466.400 ;
        RECT 1994.720 406.745 2023.070 466.400 ;
        RECT 2026.970 406.745 2055.320 466.400 ;
        RECT 2059.220 406.745 2087.570 466.400 ;
        RECT 1865.720 190.400 2087.570 406.745 ;
        RECT 1865.720 9.015 1894.070 190.400 ;
        RECT 1897.970 9.015 1926.320 190.400 ;
        RECT 1930.220 9.015 1958.570 190.400 ;
        RECT 1962.470 9.015 1990.820 190.400 ;
        RECT 1994.720 9.015 2023.070 190.400 ;
        RECT 2026.970 9.015 2055.320 190.400 ;
        RECT 2059.220 9.015 2087.570 190.400 ;
        RECT 2091.470 9.015 2119.820 3512.705 ;
        RECT 2123.720 3442.745 2152.070 3512.705 ;
        RECT 2155.970 3442.745 2184.320 3512.705 ;
        RECT 2188.220 3442.745 2216.570 3512.705 ;
        RECT 2220.470 3442.745 2248.820 3512.705 ;
        RECT 2252.720 3442.745 2281.070 3512.705 ;
        RECT 2284.970 3442.745 2313.320 3512.705 ;
        RECT 2317.220 3442.745 2345.570 3512.705 ;
        RECT 2123.720 3226.400 2345.570 3442.745 ;
        RECT 2123.720 3166.745 2152.070 3226.400 ;
        RECT 2155.970 3166.745 2184.320 3226.400 ;
        RECT 2188.220 3166.745 2216.570 3226.400 ;
        RECT 2220.470 3166.745 2248.820 3226.400 ;
        RECT 2252.720 3166.745 2281.070 3226.400 ;
        RECT 2284.970 3166.745 2313.320 3226.400 ;
        RECT 2317.220 3166.745 2345.570 3226.400 ;
        RECT 2123.720 2950.400 2345.570 3166.745 ;
        RECT 2123.720 2890.745 2152.070 2950.400 ;
        RECT 2155.970 2890.745 2184.320 2950.400 ;
        RECT 2188.220 2890.745 2216.570 2950.400 ;
        RECT 2220.470 2890.745 2248.820 2950.400 ;
        RECT 2252.720 2890.745 2281.070 2950.400 ;
        RECT 2284.970 2890.745 2313.320 2950.400 ;
        RECT 2317.220 2890.745 2345.570 2950.400 ;
        RECT 2123.720 2674.400 2345.570 2890.745 ;
        RECT 2123.720 2614.745 2152.070 2674.400 ;
        RECT 2155.970 2614.745 2184.320 2674.400 ;
        RECT 2188.220 2614.745 2216.570 2674.400 ;
        RECT 2220.470 2614.745 2248.820 2674.400 ;
        RECT 2252.720 2614.745 2281.070 2674.400 ;
        RECT 2284.970 2614.745 2313.320 2674.400 ;
        RECT 2317.220 2614.745 2345.570 2674.400 ;
        RECT 2123.720 2398.400 2345.570 2614.745 ;
        RECT 2123.720 2338.745 2152.070 2398.400 ;
        RECT 2155.970 2338.745 2184.320 2398.400 ;
        RECT 2188.220 2338.745 2216.570 2398.400 ;
        RECT 2220.470 2338.745 2248.820 2398.400 ;
        RECT 2252.720 2338.745 2281.070 2398.400 ;
        RECT 2284.970 2338.745 2313.320 2398.400 ;
        RECT 2317.220 2338.745 2345.570 2398.400 ;
        RECT 2123.720 2122.400 2345.570 2338.745 ;
        RECT 2123.720 2062.745 2152.070 2122.400 ;
        RECT 2155.970 2062.745 2184.320 2122.400 ;
        RECT 2188.220 2062.745 2216.570 2122.400 ;
        RECT 2220.470 2062.745 2248.820 2122.400 ;
        RECT 2252.720 2062.745 2281.070 2122.400 ;
        RECT 2284.970 2062.745 2313.320 2122.400 ;
        RECT 2317.220 2062.745 2345.570 2122.400 ;
        RECT 2123.720 1846.400 2345.570 2062.745 ;
        RECT 2123.720 1786.745 2152.070 1846.400 ;
        RECT 2155.970 1786.745 2184.320 1846.400 ;
        RECT 2188.220 1786.745 2216.570 1846.400 ;
        RECT 2220.470 1786.745 2248.820 1846.400 ;
        RECT 2252.720 1786.745 2281.070 1846.400 ;
        RECT 2284.970 1786.745 2313.320 1846.400 ;
        RECT 2317.220 1786.745 2345.570 1846.400 ;
        RECT 2123.720 1570.400 2345.570 1786.745 ;
        RECT 2123.720 1510.745 2152.070 1570.400 ;
        RECT 2155.970 1510.745 2184.320 1570.400 ;
        RECT 2188.220 1510.745 2216.570 1570.400 ;
        RECT 2220.470 1510.745 2248.820 1570.400 ;
        RECT 2252.720 1510.745 2281.070 1570.400 ;
        RECT 2284.970 1510.745 2313.320 1570.400 ;
        RECT 2317.220 1510.745 2345.570 1570.400 ;
        RECT 2123.720 1294.400 2345.570 1510.745 ;
        RECT 2123.720 1234.745 2152.070 1294.400 ;
        RECT 2155.970 1234.745 2184.320 1294.400 ;
        RECT 2188.220 1234.745 2216.570 1294.400 ;
        RECT 2220.470 1234.745 2248.820 1294.400 ;
        RECT 2252.720 1234.745 2281.070 1294.400 ;
        RECT 2284.970 1234.745 2313.320 1294.400 ;
        RECT 2317.220 1234.745 2345.570 1294.400 ;
        RECT 2123.720 1018.400 2345.570 1234.745 ;
        RECT 2123.720 958.745 2152.070 1018.400 ;
        RECT 2155.970 958.745 2184.320 1018.400 ;
        RECT 2188.220 958.745 2216.570 1018.400 ;
        RECT 2220.470 958.745 2248.820 1018.400 ;
        RECT 2252.720 958.745 2281.070 1018.400 ;
        RECT 2284.970 958.745 2313.320 1018.400 ;
        RECT 2317.220 958.745 2345.570 1018.400 ;
        RECT 2123.720 742.400 2345.570 958.745 ;
        RECT 2123.720 682.745 2152.070 742.400 ;
        RECT 2155.970 682.745 2184.320 742.400 ;
        RECT 2188.220 682.745 2216.570 742.400 ;
        RECT 2220.470 682.745 2248.820 742.400 ;
        RECT 2252.720 682.745 2281.070 742.400 ;
        RECT 2284.970 682.745 2313.320 742.400 ;
        RECT 2317.220 682.745 2345.570 742.400 ;
        RECT 2123.720 466.400 2345.570 682.745 ;
        RECT 2123.720 406.745 2152.070 466.400 ;
        RECT 2155.970 406.745 2184.320 466.400 ;
        RECT 2188.220 406.745 2216.570 466.400 ;
        RECT 2220.470 406.745 2248.820 466.400 ;
        RECT 2252.720 406.745 2281.070 466.400 ;
        RECT 2284.970 406.745 2313.320 466.400 ;
        RECT 2317.220 406.745 2345.570 466.400 ;
        RECT 2123.720 190.400 2345.570 406.745 ;
        RECT 2123.720 9.015 2152.070 190.400 ;
        RECT 2155.970 9.015 2184.320 190.400 ;
        RECT 2188.220 9.015 2216.570 190.400 ;
        RECT 2220.470 9.015 2248.820 190.400 ;
        RECT 2252.720 9.015 2281.070 190.400 ;
        RECT 2284.970 9.015 2313.320 190.400 ;
        RECT 2317.220 9.015 2345.570 190.400 ;
        RECT 2349.470 9.015 2377.820 3512.705 ;
        RECT 2381.720 3442.745 2410.070 3512.705 ;
        RECT 2413.970 3442.745 2442.320 3512.705 ;
        RECT 2446.220 3442.745 2474.570 3512.705 ;
        RECT 2478.470 3442.745 2506.820 3512.705 ;
        RECT 2510.720 3442.745 2539.070 3512.705 ;
        RECT 2542.970 3442.745 2571.320 3512.705 ;
        RECT 2575.220 3442.745 2603.570 3512.705 ;
        RECT 2381.720 3226.400 2603.570 3442.745 ;
        RECT 2381.720 3166.745 2410.070 3226.400 ;
        RECT 2413.970 3166.745 2442.320 3226.400 ;
        RECT 2446.220 3166.745 2474.570 3226.400 ;
        RECT 2478.470 3166.745 2506.820 3226.400 ;
        RECT 2510.720 3166.745 2539.070 3226.400 ;
        RECT 2542.970 3166.745 2571.320 3226.400 ;
        RECT 2575.220 3166.745 2603.570 3226.400 ;
        RECT 2381.720 2950.400 2603.570 3166.745 ;
        RECT 2381.720 2890.745 2410.070 2950.400 ;
        RECT 2413.970 2890.745 2442.320 2950.400 ;
        RECT 2446.220 2890.745 2474.570 2950.400 ;
        RECT 2478.470 2890.745 2506.820 2950.400 ;
        RECT 2510.720 2890.745 2539.070 2950.400 ;
        RECT 2542.970 2890.745 2571.320 2950.400 ;
        RECT 2575.220 2890.745 2603.570 2950.400 ;
        RECT 2381.720 2674.400 2603.570 2890.745 ;
        RECT 2381.720 2614.745 2410.070 2674.400 ;
        RECT 2413.970 2614.745 2442.320 2674.400 ;
        RECT 2446.220 2614.745 2474.570 2674.400 ;
        RECT 2478.470 2614.745 2506.820 2674.400 ;
        RECT 2510.720 2614.745 2539.070 2674.400 ;
        RECT 2542.970 2614.745 2571.320 2674.400 ;
        RECT 2575.220 2614.745 2603.570 2674.400 ;
        RECT 2381.720 2398.400 2603.570 2614.745 ;
        RECT 2381.720 2338.745 2410.070 2398.400 ;
        RECT 2413.970 2338.745 2442.320 2398.400 ;
        RECT 2446.220 2338.745 2474.570 2398.400 ;
        RECT 2478.470 2338.745 2506.820 2398.400 ;
        RECT 2510.720 2338.745 2539.070 2398.400 ;
        RECT 2542.970 2338.745 2571.320 2398.400 ;
        RECT 2575.220 2338.745 2603.570 2398.400 ;
        RECT 2381.720 2122.400 2603.570 2338.745 ;
        RECT 2381.720 2062.745 2410.070 2122.400 ;
        RECT 2413.970 2062.745 2442.320 2122.400 ;
        RECT 2446.220 2062.745 2474.570 2122.400 ;
        RECT 2478.470 2062.745 2506.820 2122.400 ;
        RECT 2510.720 2062.745 2539.070 2122.400 ;
        RECT 2542.970 2062.745 2571.320 2122.400 ;
        RECT 2575.220 2062.745 2603.570 2122.400 ;
        RECT 2381.720 1846.400 2603.570 2062.745 ;
        RECT 2381.720 1786.745 2410.070 1846.400 ;
        RECT 2413.970 1786.745 2442.320 1846.400 ;
        RECT 2446.220 1786.745 2474.570 1846.400 ;
        RECT 2478.470 1786.745 2506.820 1846.400 ;
        RECT 2510.720 1786.745 2539.070 1846.400 ;
        RECT 2542.970 1786.745 2571.320 1846.400 ;
        RECT 2575.220 1786.745 2603.570 1846.400 ;
        RECT 2381.720 1570.400 2603.570 1786.745 ;
        RECT 2381.720 1510.745 2410.070 1570.400 ;
        RECT 2413.970 1510.745 2442.320 1570.400 ;
        RECT 2446.220 1510.745 2474.570 1570.400 ;
        RECT 2478.470 1510.745 2506.820 1570.400 ;
        RECT 2510.720 1510.745 2539.070 1570.400 ;
        RECT 2542.970 1510.745 2571.320 1570.400 ;
        RECT 2575.220 1510.745 2603.570 1570.400 ;
        RECT 2381.720 1294.400 2603.570 1510.745 ;
        RECT 2381.720 1234.745 2410.070 1294.400 ;
        RECT 2413.970 1234.745 2442.320 1294.400 ;
        RECT 2446.220 1234.745 2474.570 1294.400 ;
        RECT 2478.470 1234.745 2506.820 1294.400 ;
        RECT 2510.720 1234.745 2539.070 1294.400 ;
        RECT 2542.970 1234.745 2571.320 1294.400 ;
        RECT 2575.220 1234.745 2603.570 1294.400 ;
        RECT 2381.720 1018.400 2603.570 1234.745 ;
        RECT 2381.720 958.745 2410.070 1018.400 ;
        RECT 2413.970 958.745 2442.320 1018.400 ;
        RECT 2446.220 958.745 2474.570 1018.400 ;
        RECT 2478.470 958.745 2506.820 1018.400 ;
        RECT 2510.720 958.745 2539.070 1018.400 ;
        RECT 2542.970 958.745 2571.320 1018.400 ;
        RECT 2575.220 958.745 2603.570 1018.400 ;
        RECT 2381.720 742.400 2603.570 958.745 ;
        RECT 2381.720 682.745 2410.070 742.400 ;
        RECT 2413.970 682.745 2442.320 742.400 ;
        RECT 2446.220 682.745 2474.570 742.400 ;
        RECT 2478.470 682.745 2506.820 742.400 ;
        RECT 2510.720 682.745 2539.070 742.400 ;
        RECT 2542.970 682.745 2571.320 742.400 ;
        RECT 2575.220 682.745 2603.570 742.400 ;
        RECT 2381.720 466.400 2603.570 682.745 ;
        RECT 2381.720 406.745 2410.070 466.400 ;
        RECT 2413.970 406.745 2442.320 466.400 ;
        RECT 2446.220 406.745 2474.570 466.400 ;
        RECT 2478.470 406.745 2506.820 466.400 ;
        RECT 2510.720 406.745 2539.070 466.400 ;
        RECT 2542.970 406.745 2571.320 466.400 ;
        RECT 2575.220 406.745 2603.570 466.400 ;
        RECT 2381.720 190.400 2603.570 406.745 ;
        RECT 2381.720 9.015 2410.070 190.400 ;
        RECT 2413.970 9.015 2442.320 190.400 ;
        RECT 2446.220 9.015 2474.570 190.400 ;
        RECT 2478.470 9.015 2506.820 190.400 ;
        RECT 2510.720 9.015 2539.070 190.400 ;
        RECT 2542.970 9.015 2571.320 190.400 ;
        RECT 2575.220 9.015 2603.570 190.400 ;
        RECT 2607.470 9.015 2635.820 3512.705 ;
        RECT 2639.720 3442.745 2668.070 3512.705 ;
        RECT 2671.970 3442.745 2700.320 3512.705 ;
        RECT 2704.220 3442.745 2732.570 3512.705 ;
        RECT 2736.470 3442.745 2764.820 3512.705 ;
        RECT 2768.720 3442.745 2797.070 3512.705 ;
        RECT 2800.970 3442.745 2829.320 3512.705 ;
        RECT 2833.220 3442.745 2861.570 3512.705 ;
        RECT 2639.720 3226.400 2861.570 3442.745 ;
        RECT 2639.720 3166.745 2668.070 3226.400 ;
        RECT 2671.970 3166.745 2700.320 3226.400 ;
        RECT 2704.220 3166.745 2732.570 3226.400 ;
        RECT 2736.470 3166.745 2764.820 3226.400 ;
        RECT 2768.720 3166.745 2797.070 3226.400 ;
        RECT 2800.970 3166.745 2829.320 3226.400 ;
        RECT 2833.220 3166.745 2861.570 3226.400 ;
        RECT 2639.720 2950.400 2861.570 3166.745 ;
        RECT 2639.720 2890.745 2668.070 2950.400 ;
        RECT 2671.970 2890.745 2700.320 2950.400 ;
        RECT 2704.220 2890.745 2732.570 2950.400 ;
        RECT 2736.470 2890.745 2764.820 2950.400 ;
        RECT 2768.720 2890.745 2797.070 2950.400 ;
        RECT 2800.970 2890.745 2829.320 2950.400 ;
        RECT 2833.220 2890.745 2861.570 2950.400 ;
        RECT 2639.720 2674.400 2861.570 2890.745 ;
        RECT 2639.720 2614.745 2668.070 2674.400 ;
        RECT 2671.970 2614.745 2700.320 2674.400 ;
        RECT 2704.220 2614.745 2732.570 2674.400 ;
        RECT 2736.470 2614.745 2764.820 2674.400 ;
        RECT 2768.720 2614.745 2797.070 2674.400 ;
        RECT 2800.970 2614.745 2829.320 2674.400 ;
        RECT 2833.220 2614.745 2861.570 2674.400 ;
        RECT 2639.720 2398.400 2861.570 2614.745 ;
        RECT 2639.720 2338.745 2668.070 2398.400 ;
        RECT 2671.970 2338.745 2700.320 2398.400 ;
        RECT 2704.220 2338.745 2732.570 2398.400 ;
        RECT 2736.470 2338.745 2764.820 2398.400 ;
        RECT 2768.720 2338.745 2797.070 2398.400 ;
        RECT 2800.970 2338.745 2829.320 2398.400 ;
        RECT 2833.220 2338.745 2861.570 2398.400 ;
        RECT 2639.720 2122.400 2861.570 2338.745 ;
        RECT 2639.720 2062.745 2668.070 2122.400 ;
        RECT 2671.970 2062.745 2700.320 2122.400 ;
        RECT 2704.220 2062.745 2732.570 2122.400 ;
        RECT 2736.470 2062.745 2764.820 2122.400 ;
        RECT 2768.720 2062.745 2797.070 2122.400 ;
        RECT 2800.970 2062.745 2829.320 2122.400 ;
        RECT 2833.220 2062.745 2861.570 2122.400 ;
        RECT 2639.720 1846.400 2861.570 2062.745 ;
        RECT 2639.720 1786.745 2668.070 1846.400 ;
        RECT 2671.970 1786.745 2700.320 1846.400 ;
        RECT 2704.220 1786.745 2732.570 1846.400 ;
        RECT 2736.470 1786.745 2764.820 1846.400 ;
        RECT 2768.720 1786.745 2797.070 1846.400 ;
        RECT 2800.970 1786.745 2829.320 1846.400 ;
        RECT 2833.220 1786.745 2861.570 1846.400 ;
        RECT 2639.720 1570.400 2861.570 1786.745 ;
        RECT 2639.720 1510.745 2668.070 1570.400 ;
        RECT 2671.970 1510.745 2700.320 1570.400 ;
        RECT 2704.220 1510.745 2732.570 1570.400 ;
        RECT 2736.470 1510.745 2764.820 1570.400 ;
        RECT 2768.720 1510.745 2797.070 1570.400 ;
        RECT 2800.970 1510.745 2829.320 1570.400 ;
        RECT 2833.220 1510.745 2861.570 1570.400 ;
        RECT 2639.720 1294.400 2861.570 1510.745 ;
        RECT 2639.720 1234.745 2668.070 1294.400 ;
        RECT 2671.970 1234.745 2700.320 1294.400 ;
        RECT 2704.220 1234.745 2732.570 1294.400 ;
        RECT 2736.470 1234.745 2764.820 1294.400 ;
        RECT 2768.720 1234.745 2797.070 1294.400 ;
        RECT 2800.970 1234.745 2829.320 1294.400 ;
        RECT 2833.220 1234.745 2861.570 1294.400 ;
        RECT 2639.720 1018.400 2861.570 1234.745 ;
        RECT 2639.720 958.745 2668.070 1018.400 ;
        RECT 2671.970 958.745 2700.320 1018.400 ;
        RECT 2704.220 958.745 2732.570 1018.400 ;
        RECT 2736.470 958.745 2764.820 1018.400 ;
        RECT 2768.720 958.745 2797.070 1018.400 ;
        RECT 2800.970 958.745 2829.320 1018.400 ;
        RECT 2833.220 958.745 2861.570 1018.400 ;
        RECT 2639.720 742.400 2861.570 958.745 ;
        RECT 2639.720 682.745 2668.070 742.400 ;
        RECT 2671.970 682.745 2700.320 742.400 ;
        RECT 2704.220 682.745 2732.570 742.400 ;
        RECT 2736.470 682.745 2764.820 742.400 ;
        RECT 2768.720 682.745 2797.070 742.400 ;
        RECT 2800.970 682.745 2829.320 742.400 ;
        RECT 2833.220 682.745 2861.570 742.400 ;
        RECT 2639.720 466.400 2861.570 682.745 ;
        RECT 2639.720 406.745 2668.070 466.400 ;
        RECT 2671.970 406.745 2700.320 466.400 ;
        RECT 2704.220 406.745 2732.570 466.400 ;
        RECT 2736.470 406.745 2764.820 466.400 ;
        RECT 2768.720 406.745 2797.070 466.400 ;
        RECT 2800.970 406.745 2829.320 466.400 ;
        RECT 2833.220 406.745 2861.570 466.400 ;
        RECT 2639.720 190.400 2861.570 406.745 ;
        RECT 2639.720 9.015 2668.070 190.400 ;
        RECT 2671.970 9.015 2700.320 190.400 ;
        RECT 2704.220 9.015 2732.570 190.400 ;
        RECT 2736.470 9.015 2764.820 190.400 ;
        RECT 2768.720 9.015 2797.070 190.400 ;
        RECT 2800.970 9.015 2829.320 190.400 ;
        RECT 2833.220 9.015 2861.570 190.400 ;
        RECT 2865.470 9.015 2893.820 3512.705 ;
        RECT 2897.720 9.015 2911.505 3512.705 ;
      LAYER met5 ;
        RECT 18.980 3452.280 2869.820 3460.300 ;
        RECT 18.980 3435.030 2869.820 3445.980 ;
        RECT 18.980 3417.780 2869.820 3428.730 ;
        RECT 18.980 3400.530 2869.820 3411.480 ;
        RECT 18.980 3383.280 2869.820 3394.230 ;
        RECT 18.980 3366.030 2869.820 3376.980 ;
        RECT 18.980 3348.780 2869.820 3359.730 ;
        RECT 18.980 3331.530 2869.820 3342.480 ;
        RECT 18.980 3314.280 2869.820 3325.230 ;
        RECT 18.980 3297.030 2869.820 3307.980 ;
        RECT 18.980 3279.780 2869.820 3290.730 ;
        RECT 18.980 3262.530 2869.820 3273.480 ;
        RECT 18.980 3245.280 2869.820 3256.230 ;
        RECT 18.980 3228.030 2869.820 3238.980 ;
        RECT 18.980 3210.780 2869.820 3221.730 ;
        RECT 18.980 3193.530 2869.820 3204.480 ;
        RECT 18.980 3176.280 2869.820 3187.230 ;
        RECT 18.980 3159.030 2869.820 3169.980 ;
        RECT 18.980 3141.780 2869.820 3152.730 ;
        RECT 18.980 3124.530 2869.820 3135.480 ;
        RECT 18.980 3107.280 2869.820 3118.230 ;
        RECT 18.980 3090.030 2869.820 3100.980 ;
        RECT 18.980 3072.780 2869.820 3083.730 ;
        RECT 18.980 3055.530 2869.820 3066.480 ;
        RECT 18.980 3038.280 2869.820 3049.230 ;
        RECT 18.980 3021.030 2869.820 3031.980 ;
        RECT 18.980 3003.780 2869.820 3014.730 ;
        RECT 18.980 2986.530 2869.820 2997.480 ;
        RECT 18.980 2969.280 2869.820 2980.230 ;
        RECT 18.980 2952.030 2869.820 2962.980 ;
        RECT 18.980 2934.780 2869.820 2945.730 ;
        RECT 18.980 2917.530 2869.820 2928.480 ;
        RECT 18.980 2900.280 2869.820 2911.230 ;
        RECT 18.980 2883.030 2869.820 2893.980 ;
        RECT 18.980 2865.780 2869.820 2876.730 ;
        RECT 18.980 2848.530 2869.820 2859.480 ;
        RECT 18.980 2831.280 2869.820 2842.230 ;
        RECT 18.980 2814.030 2869.820 2824.980 ;
        RECT 18.980 2796.780 2869.820 2807.730 ;
        RECT 18.980 2779.530 2869.820 2790.480 ;
        RECT 18.980 2762.280 2869.820 2773.230 ;
        RECT 18.980 2745.030 2869.820 2755.980 ;
        RECT 18.980 2727.780 2869.820 2738.730 ;
        RECT 18.980 2710.530 2869.820 2721.480 ;
        RECT 18.980 2693.280 2869.820 2704.230 ;
        RECT 18.980 2676.030 2869.820 2686.980 ;
        RECT 18.980 2658.780 2869.820 2669.730 ;
        RECT 18.980 2641.530 2869.820 2652.480 ;
        RECT 18.980 2624.280 2869.820 2635.230 ;
        RECT 18.980 2607.030 2869.820 2617.980 ;
        RECT 18.980 2589.780 2869.820 2600.730 ;
        RECT 18.980 2572.530 2869.820 2583.480 ;
        RECT 18.980 2555.280 2869.820 2566.230 ;
        RECT 18.980 2538.030 2869.820 2548.980 ;
        RECT 18.980 2520.780 2869.820 2531.730 ;
        RECT 18.980 2503.530 2869.820 2514.480 ;
        RECT 18.980 2486.280 2869.820 2497.230 ;
        RECT 18.980 2469.030 2869.820 2479.980 ;
        RECT 18.980 2451.780 2869.820 2462.730 ;
        RECT 18.980 2434.530 2869.820 2445.480 ;
        RECT 18.980 2417.280 2869.820 2428.230 ;
        RECT 18.980 2400.030 2869.820 2410.980 ;
        RECT 18.980 2382.780 2869.820 2393.730 ;
        RECT 18.980 2365.530 2869.820 2376.480 ;
        RECT 18.980 2348.280 2869.820 2359.230 ;
        RECT 18.980 2331.030 2869.820 2341.980 ;
        RECT 18.980 2313.780 2869.820 2324.730 ;
        RECT 18.980 2296.530 2869.820 2307.480 ;
        RECT 18.980 2279.280 2869.820 2290.230 ;
        RECT 18.980 2262.030 2869.820 2272.980 ;
        RECT 18.980 2244.780 2869.820 2255.730 ;
        RECT 18.980 2227.530 2869.820 2238.480 ;
        RECT 18.980 2210.280 2869.820 2221.230 ;
        RECT 18.980 2193.030 2869.820 2203.980 ;
        RECT 18.980 2175.780 2869.820 2186.730 ;
        RECT 18.980 2158.530 2869.820 2169.480 ;
        RECT 18.980 2141.280 2869.820 2152.230 ;
        RECT 18.980 2124.030 2869.820 2134.980 ;
        RECT 18.980 2106.780 2869.820 2117.730 ;
        RECT 18.980 2089.530 2869.820 2100.480 ;
        RECT 18.980 2072.280 2869.820 2083.230 ;
        RECT 18.980 2055.030 2869.820 2065.980 ;
        RECT 18.980 2037.780 2869.820 2048.730 ;
        RECT 18.980 2020.530 2869.820 2031.480 ;
        RECT 18.980 2003.280 2869.820 2014.230 ;
        RECT 18.980 1986.030 2869.820 1996.980 ;
        RECT 18.980 1968.780 2869.820 1979.730 ;
        RECT 18.980 1951.530 2869.820 1962.480 ;
        RECT 18.980 1934.280 2869.820 1945.230 ;
        RECT 18.980 1917.030 2869.820 1927.980 ;
        RECT 18.980 1899.780 2869.820 1910.730 ;
        RECT 18.980 1882.530 2869.820 1893.480 ;
        RECT 18.980 1865.280 2869.820 1876.230 ;
        RECT 18.980 1848.030 2869.820 1858.980 ;
        RECT 18.980 1830.780 2869.820 1841.730 ;
        RECT 18.980 1813.530 2869.820 1824.480 ;
        RECT 18.980 1796.280 2869.820 1807.230 ;
        RECT 18.980 1779.030 2869.820 1789.980 ;
        RECT 18.980 1761.780 2869.820 1772.730 ;
        RECT 18.980 1744.530 2869.820 1755.480 ;
        RECT 18.980 1727.280 2869.820 1738.230 ;
        RECT 18.980 1710.030 2869.820 1720.980 ;
        RECT 18.980 1692.780 2869.820 1703.730 ;
        RECT 18.980 1675.530 2869.820 1686.480 ;
        RECT 18.980 1658.280 2869.820 1669.230 ;
        RECT 18.980 1641.030 2869.820 1651.980 ;
        RECT 18.980 1623.780 2869.820 1634.730 ;
        RECT 18.980 1606.530 2869.820 1617.480 ;
        RECT 18.980 1589.280 2869.820 1600.230 ;
        RECT 18.980 1572.030 2869.820 1582.980 ;
        RECT 18.980 1554.780 2869.820 1565.730 ;
        RECT 18.980 1537.530 2869.820 1548.480 ;
        RECT 18.980 1520.280 2869.820 1531.230 ;
        RECT 18.980 1503.030 2869.820 1513.980 ;
        RECT 18.980 1485.780 2869.820 1496.730 ;
        RECT 18.980 1468.530 2869.820 1479.480 ;
        RECT 18.980 1451.280 2869.820 1462.230 ;
        RECT 18.980 1434.030 2869.820 1444.980 ;
        RECT 18.980 1416.780 2869.820 1427.730 ;
        RECT 18.980 1399.530 2869.820 1410.480 ;
        RECT 18.980 1382.280 2869.820 1393.230 ;
        RECT 18.980 1365.030 2869.820 1375.980 ;
        RECT 18.980 1347.780 2869.820 1358.730 ;
        RECT 18.980 1330.530 2869.820 1341.480 ;
        RECT 18.980 1313.280 2869.820 1324.230 ;
        RECT 18.980 1296.030 2869.820 1306.980 ;
        RECT 18.980 1278.780 2869.820 1289.730 ;
        RECT 18.980 1261.530 2869.820 1272.480 ;
        RECT 18.980 1244.280 2869.820 1255.230 ;
        RECT 18.980 1227.030 2869.820 1237.980 ;
        RECT 18.980 1209.780 2869.820 1220.730 ;
        RECT 18.980 1192.530 2869.820 1203.480 ;
        RECT 18.980 1175.280 2869.820 1186.230 ;
        RECT 18.980 1158.030 2869.820 1168.980 ;
        RECT 18.980 1140.780 2869.820 1151.730 ;
        RECT 18.980 1123.530 2869.820 1134.480 ;
        RECT 18.980 1106.280 2869.820 1117.230 ;
        RECT 18.980 1089.030 2869.820 1099.980 ;
        RECT 18.980 1071.780 2869.820 1082.730 ;
        RECT 18.980 1054.530 2869.820 1065.480 ;
        RECT 18.980 1037.280 2869.820 1048.230 ;
        RECT 18.980 1020.030 2869.820 1030.980 ;
        RECT 18.980 1002.780 2869.820 1013.730 ;
        RECT 18.980 985.530 2869.820 996.480 ;
        RECT 18.980 968.280 2869.820 979.230 ;
        RECT 18.980 951.030 2869.820 961.980 ;
        RECT 18.980 933.780 2869.820 944.730 ;
        RECT 18.980 916.530 2869.820 927.480 ;
        RECT 18.980 899.280 2869.820 910.230 ;
        RECT 18.980 882.030 2869.820 892.980 ;
        RECT 18.980 864.780 2869.820 875.730 ;
        RECT 18.980 847.530 2869.820 858.480 ;
        RECT 18.980 830.280 2869.820 841.230 ;
        RECT 18.980 813.030 2869.820 823.980 ;
        RECT 18.980 795.780 2869.820 806.730 ;
        RECT 18.980 778.530 2869.820 789.480 ;
        RECT 18.980 761.280 2869.820 772.230 ;
        RECT 18.980 744.030 2869.820 754.980 ;
        RECT 18.980 726.780 2869.820 737.730 ;
        RECT 18.980 709.530 2869.820 720.480 ;
        RECT 18.980 692.280 2869.820 703.230 ;
        RECT 18.980 675.030 2869.820 685.980 ;
        RECT 18.980 657.780 2869.820 668.730 ;
        RECT 18.980 640.530 2869.820 651.480 ;
        RECT 18.980 623.280 2869.820 634.230 ;
        RECT 18.980 606.030 2869.820 616.980 ;
        RECT 18.980 588.780 2869.820 599.730 ;
        RECT 18.980 571.530 2869.820 582.480 ;
        RECT 18.980 554.280 2869.820 565.230 ;
        RECT 18.980 537.030 2869.820 547.980 ;
        RECT 18.980 519.780 2869.820 530.730 ;
        RECT 18.980 502.530 2869.820 513.480 ;
        RECT 18.980 485.280 2869.820 496.230 ;
        RECT 18.980 468.030 2869.820 478.980 ;
        RECT 18.980 450.780 2869.820 461.730 ;
        RECT 18.980 433.530 2869.820 444.480 ;
        RECT 18.980 416.280 2869.820 427.230 ;
        RECT 18.980 399.030 2869.820 409.980 ;
        RECT 18.980 381.780 2869.820 392.730 ;
        RECT 18.980 364.530 2869.820 375.480 ;
        RECT 18.980 347.280 2869.820 358.230 ;
        RECT 18.980 330.030 2869.820 340.980 ;
        RECT 18.980 312.780 2869.820 323.730 ;
        RECT 18.980 295.530 2869.820 306.480 ;
        RECT 18.980 278.280 2869.820 289.230 ;
        RECT 18.980 261.030 2869.820 271.980 ;
        RECT 18.980 243.780 2869.820 254.730 ;
        RECT 18.980 226.530 2869.820 237.480 ;
        RECT 18.980 209.280 2869.820 220.230 ;
        RECT 18.980 192.030 2869.820 202.980 ;
        RECT 18.980 174.780 2869.820 185.730 ;
        RECT 18.980 157.530 2869.820 168.480 ;
        RECT 18.980 140.280 2869.820 151.230 ;
        RECT 18.980 123.030 2869.820 133.980 ;
        RECT 18.980 105.780 2869.820 116.730 ;
        RECT 18.980 88.530 2869.820 99.480 ;
        RECT 18.980 71.280 2869.820 82.230 ;
        RECT 18.980 54.030 2869.820 64.980 ;
        RECT 18.980 21.300 2869.820 47.730 ;
  END
END user_project_wrapper
END LIBRARY

